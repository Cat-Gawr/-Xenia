library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package pixelNum_pkg is
type pixArray is array (0 to 47, 0 to 47) of std_logic_vector(23 downto 0);
constant pix0: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);

constant pix1: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);

constant pix2: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);


constant pix3: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);


constant pix4: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);


constant pix5: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);


constant pix6: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);


constant pix7: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);

constant pix8: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);

constant pix9: pixArray := (
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"E38029", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"5C2814", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000"),
    (X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000", X"000000")
);


end pixelNum_pkg;
