library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package endgame_pkg is
    type overArray is array (0 to 67, 0 to 87) of std_logic_vector(23 downto 0);
    type winArray is array (0 to 11, 0 to 59) of std_logic_vector(23 downto 0);
    type LOGOArray is array (0 to 180, 0 to 267) of std_logic_vector(23 downto 0);

    constant over: overArray := (
        (X"F9FFE6", X"F8FFEB", X"F4FFF2", X"F2FBFA", X"DFE8F3", X"5E697A", X"586577", X"5E6A7F", X"5A6779", X"5A6777", X"5A6777", X"596676", X"586575", X"586374", X"5A6274", X"5B6176", X"5F627A", X"575669", X"929196", X"FBF7F6", X"FEF8F5", X"FFFBFB", X"FEF4FC", X"FFF7FF", X"FDFAFF", X"B9B9C4", X"51576C", X"575C75", X"5E5C78", X"645974", X"6E566A", X"6C566E", X"5E5B7C", X"565F7C", X"56626E", X"566366", X"586762", X"54625F", X"4E5B5F", X"AFB2BA", X"FFF9FF", X"FFF1FF", X"FFF0FF", X"FBEBFF", X"747187", X"61637B", X"595C84", X"5E6291", X"5E638F", X"595F7F", X"6C747A", X"EFF7ED", X"F6FEE9", X"FAFFEB", X"FFFFFF", X"FFFFFB", X"F6F4F2", X"FEFCFD", X"FAF7FA", X"FCF8FF", X"77757F", X"646471", X"727484", X"656B7B", X"576072", X"55606E", X"606A72", X"E1EBF1", X"F2FDFF", X"8C969E", X"4D5866", X"5A6276", X"615F79", X"635F79", X"606079", X"5D6279", X"586479", X"536779", X"506879", X"55657D", X"605E83", X"635D7F", X"606175", X"5E646B", X"525C56", X"B1BEB3", X"F5FFF7", X"EBF9ED"),
        (X"F1FAE2", X"F8FFEF", X"FFFFFE", X"FFFFFF", X"D5DBE0", X"131C20", X"0F1719", X"131A17", X"131814", X"131912", X"131912", X"121711", X"111610", X"0F150F", X"11140F", X"131311", X"161616", X"020000", X"66625F", X"FFFEF9", X"FFFFFF", X"FFFDFF", X"FFF7FF", X"FFFBFF", X"FEFBFF", X"97999B", X"000006", X"18171F", X"170F17", X"1C0E11", X"230C0B", X"1F0D0D", X"161019", X"111317", X"11150D", X"111605", X"111702", X"131907", X"0A0E06", X"949293", X"FFFFFF", X"FFF9FF", X"FFF5FF", X"FEF2FF", X"1D171E", X"141316", X"110F1E", X"121124", X"16182A", X"010612", X"2B3232", X"F2F8F0", X"F9FFF3", X"F2F6E9", X"FAFDF5", X"FFFFFB", X"FEFCFB", X"FCFAFA", X"FFFFFF", X"FFFFFF", X"332F2A", X"15150A", X"13140D", X"171815", X"111411", X"121715", X"212526", X"ECF0F3", X"FCFFFF", X"6A6F6F", X"000200", X"161817", X"150D12", X"150D14", X"130E14", X"101014", X"0C1214", X"081414", X"051514", X"081316", X"120E1A", X"150D16", X"12100E", X"101208", X"000400", X"8C9584", X"F6FFF5", X"FBFFFC"),
        (X"F6FAF0", X"FDFFF9", X"DADCDE", X"A4A4A6", X"9C9B97", X"696A57", X"6F714C", X"7A7849", X"766E3D", X"786E3B", X"786E3B", X"776D3A", X"766C38", X"746B37", X"746B37", X"736B39", X"746B3E", X"69613D", X"837C65", X"ACA298", X"B4AAAD", X"FFFDFF", X"FFFBFF", X"C4BEC7", X"ABACA7", X"8C8C7E", X"716953", X"726547", X"7D6A45", X"7E6A41", X"7D6B3F", X"7B6B41", X"796B45", X"796C43", X"796D3B", X"796E39", X"716533", X"716439", X"6F5F42", X"958777", X"AAA4A1", X"A29FA7", X"A29EAD", X"ABA4A9", X"6F654D", X"796D46", X"7B6F4A", X"766C49", X"71704C", X"747658", X"717164", X"A5A6A1", X"ACACAE", X"E7E9ED", X"F2F4F3", X"F1F1EF", X"FDFDFB", X"E6E3E6", X"A39CA8", X"AEA7A5", X"706E44", X"716F34", X"686232", X"716B3F", X"6D663B", X"706748", X"6E6558", X"A09894", X"ACA39F", X"837A6D", X"726A4B", X"7D7149", X"796844", X"796747", X"776847", X"766947", X"746A47", X"716B47", X"6F6C47", X"716B47", X"746A47", X"766944", X"766B3E", X"726C3E", X"646139", X"919375", X"ABB5A4", X"B4BFB4"),
        (X"FFFFFF", X"FFFFFF", X"9F9A9E", X"160D09", X"453D26", X"E6DDB3", X"F3EDA6", X"E4D986", X"F8E38F", X"FBE28D", X"FBE28D", X"FAE18C", X"F8DF8B", X"F6DF89", X"F6DF89", X"F4E08B", X"E4D483", X"F9EBA9", X"AD9F74", X"120600", X"342624", X"EFE5ED", X"FFFBFF", X"5D585A", X"020300", X"726F49", X"FDEFBB", X"F4DC9C", X"F5DA8F", X"F5DB8B", X"F0DD8D", X"F0DD8F", X"F3DB91", X"F6DA8D", X"F6DB87", X"F6DB87", X"FFE79A", X"FCDE9B", X"FFE5B2", X"745C39", X"141000", X"131814", X"1C2025", X"2A261E", X"DCCB9A", X"F2DB93", X"F9E396", X"EEDE8F", X"E0D889", X"F2ECAC", X"CCC5A7", X"2D2420", X"1E1823", X"B7B5C1", X"FFFFFF", X"F8FAF7", X"F5F8F7", X"CCC9CD", X"160D1A", X"1F160B", X"BEB977", X"F1EC90", X"F0E492", X"EFE093", X"F0DE92", X"EFDEA2", X"E5D5B8", X"332318", X"150400", X"A59377", X"FFECB1", X"F6E098", X"F9E09B", X"F9E09B", X"F9E09B", X"F9E09B", X"F8E19B", X"F8E19B", X"F6E29B", X"F6E29B", X"F8E19B", X"F8E199", X"F9E195", X"F6E29B", X"FFF3BB", X"7C744E", X"101304", X"4A524D"),
        (X"DFD8E8", X"E8DFE9", X"A49998", X"32230F", X"6F5D31", X"E6D48D", X"EAD574", X"F0D769", X"F0D062", X"EFCA5D", X"F1CC60", X"F7D266", X"F4CF63", X"FDDB6E", X"EECC5F", X"F4D368", X"ECD568", X"EEDB7D", X"C1AE6E", X"44310A", X"544437", X"DCD0D2", X"F8F0F7", X"706A63", X"373206", X"8E8540", X"E7D37F", X"F3D878", X"F7D66D", X"E9CB5C", X"F0D769", X"E3C95E", X"F0CC69", X"EDC460", X"EDC55A", X"F3CB60", X"F4CB67", X"F3C86E", X"FFDE92", X"9E7F43", X"413C13", X"343C25", X"232A26", X"3F3B28", X"E3C987", X"F5D273", X"EED169", X"EFD86A", X"D8C656", X"F2E389", X"D8C698", X"3B2B1E", X"271D25", X"C9C4D1", X"FCFFFE", X"FFFFFF", X"F2F4F5", X"D1CED3", X"2F242F", X"332613", X"CEC370", X"EBDE6E", X"E8D366", X"EFD56C", X"EFD26C", X"EFD482", X"DBC49A", X"4B3823", X"261300", X"A79166", X"FADE8D", X"F1D16C", X"F0D370", X"F0D372", X"F2D272", X"F4D172", X"F2D070", X"F0CB6D", X"EDC869", X"ECC768", X"EEC96B", X"F0CC6B", X"F4CB69", X"F0CB71", X"F6D895", X"8C7A50", X"221C15", X"53565E"),
        (X"5E546C", X"251823", X"7B6B5E", X"E0CDA6", X"E1CB85", X"EED174", X"F1D161", X"FED961", X"FCD15D", X"FFD363", X"FFD262", X"FDD05F", X"FDD05F", X"FFD464", X"FBCD5D", X"FBD261", X"F4D25E", X"F7DB71", X"F6DD8A", X"E3CE96", X"C9B99A", X"3C3024", X"2A2524", X"A59F8C", X"DED48F", X"E4D571", X"F2DA6E", X"EDD05D", X"F6D65B", X"F3D152", X"F8D657", X"F5D056", X"FFD468", X"FFD56C", X"FFD361", X"FACB57", X"FFD05F", X"FFD169", X"FFD175", X"EAC574", X"DED493", X"959A6E", X"111B0A", X"323013", X"E8C97D", X"FBD169", X"F1D25F", X"F3D960", X"E8CF51", X"F3D970", X"D1B97D", X"3F2A11", X"281B18", X"C1BCC0", X"F7FDF6", X"F3FBF4", X"FDFFFF", X"D8D4DC", X"1F1317", X"39290F", X"D3C16E", X"F2DB6A", X"F0D15C", X"F7D35D", X"F6D25E", X"F4D476", X"DCC591", X"4B3A1B", X"261400", X"A9925E", X"FFDE80", X"F6D160", X"F4D463", X"F4D463", X"F5D363", X"F7D062", X"F9CF62", X"FED065", X"FFD469", X"FFD36B", X"FFD06A", X"FFCC68", X"FFCC63", X"FFCA6E", X"FFDC97", X"90724C", X"1E1214", X"575469"),
        (X"574C69", X"160912", X"806E50", X"FFECAB", X"F2D677", X"F1CC5E", X"FDD25F", X"F9C958", X"FFCF67", X"FFCD6A", X"FFCF6C", X"FFD471", X"FFCD6A", X"FCCB67", X"FFD471", X"FFD972", X"FFD568", X"F4D166", X"F0D274", X"EFDA8B", X"DDCF98", X"3C3312", X"1E1B11", X"AEA888", X"F8E585", X"ECD355", X"EBD458", X"EFD65A", X"F1D357", X"FDD759", X"FECF4D", X"FFD359", X"FFD878", X"FFCE73", X"FECA63", X"FFCD5C", X"FFD360", X"FFCF61", X"FFCC64", X"FFDB7B", X"F4E386", X"A4A25E", X"131700", X"3C3618", X"EBC77D", X"FDCF6D", X"F0D169", X"F1D86A", X"EBCA53", X"FBD86F", X"D6B671", X"3D2300", X"281807", X"BFBCB1", X"FFFFFC", X"F2FCF2", X"F9FDFF", X"D1CDD5", X"241914", X"251100", X"D8BC78", X"F8D578", X"F8CE63", X"FDD05D", X"F9D05E", X"F5D577", X"DAC891", X"483C17", X"231700", X"A6945C", X"FFDE80", X"F6D160", X"F4D463", X"F2D563", X"F5D363", X"F7D062", X"FCCE62", X"FFCD63", X"FFD068", X"FFD16F", X"FFD176", X"FFCF76", X"FFCD70", X"FFCD7A", X"FFD297", X"9B6F55", X"240F1F", X"51496B"),
        (X"5D526F", X"14070E", X"857349", X"F8E092", X"F2D266", X"FFD760", X"F3C653", X"FCC95F", X"FFD774", X"D9A147", X"C27D2D", X"CA8236", X"BB7626", X"CE8C39", X"FFC36B", X"FFC96A", X"FFD06A", X"FCD46B", X"F6CF6C", X"E9C977", X"D6C287", X"3F330E", X"2C2314", X"AA9C76", X"F4D76F", X"F2D14B", X"E7CE50", X"F0D85F", X"F9DB61", X"F6CA52", X"D2931F", X"CA801C", X"C87B31", X"BC742D", X"D5963C", X"FFCC63", X"FECE5C", X"F6CB58", X"FDD163", X"F4CF65", X"F6E07A", X"ADA357", X"212106", X"342B0E", X"EBC77D", X"FBD06D", X"F0D169", X"F3D76A", X"FFD966", X"F6CF63", X"F9D783", X"B89D60", X"C7B78C", X"736D4F", X"51523B", X"5F6357", X"575958", X"6D6964", X"B4A789", X"B59D6A", X"DBBC72", X"F9D176", X"F9CE5F", X"FDD05B", X"F8CF5B", X"F5D673", X"DCC88D", X"473B14", X"211700", X"A4945E", X"FFDE80", X"F6D160", X"F2D55F", X"F2D561", X"F7D263", X"FDCE66", X"CB902D", X"CE892C", X"CF822A", X"CE7E2C", X"CD7E34", X"D17D37", X"D77B31", X"D47B39", X"CA8050", X"7C4936", X"1E091C", X"4B446B"),
        (X"554C66", X"1E1214", X"847244", X"F7DE8B", X"F5D467", X"F9D45F", X"F9D267", X"FBD06B", X"FFD270", X"DB9848", X"BD5526", X"CB5934", X"BF5826", X"BE5F22", X"FFAB60", X"FFD079", X"FFD775", X"FFD975", X"FFD57B", X"FFD38D", X"E5C398", X"462C15", X"251003", X"BCA27D", X"FED775", X"F5CE53", X"F0D65F", X"F2DA67", X"F4D25E", X"FDCA60", X"CA7826", X"C25A1D", X"CB542F", X"C05129", X"C8732E", X"FFC268", X"F8CE61", X"F2D35E", X"F1D45E", X"EFD464", X"F5DE7B", X"B7A764", X"231809", X"392C19", X"E6CA7B", X"F6D465", X"F3D15F", X"F8D461", X"FCD462", X"F9CF62", X"F6D36B", X"EED479", X"F2E099", X"4C400D", X"170B00", X"261D0E", X"171305", X"3F3916", X"F5E39E", X"EBD175", X"F5D072", X"F9D267", X"F6D356", X"F7D553", X"F3D156", X"F7D772", X"E0C988", X"493911", X"211600", X"A39366", X"FFDD86", X"F6D160", X"EFD85B", X"F0D75B", X"FAD161", X"FFCA68", X"CC7C2A", X"BB5914", X"C65519", X"C85621", X"C15A27", X"C05829", X"C9522A", X"C3522D", X"BC6241", X"773C29", X"271723", X"4B506C"),
        (X"534D64", X"1D1412", X"847342", X"F9DD89", X"F6D467", X"F9D45F", X"F8D269", X"F9D16D", X"FFD26E", X"DE9748", X"C3502E", X"D5523E", X"CA5230", X"CA5F2C", X"EA8746", X"F39E52", X"E09E47", X"DE9E49", X"E49A4D", X"E0995F", X"C19174", X"4E2D21", X"321B10", X"BAA37D", X"FCD779", X"F4CF55", X"EFD663", X"F1DA69", X"F4D260", X"FFC766", X"CF7332", X"C8542E", X"DA5741", X"D0553A", X"D3783E", X"FFCB75", X"F7D064", X"EFD55E", X"EED65E", X"ECD564", X"F5DE7D", X"BBA566", X"25160E", X"3A2A1D", X"E3CC7B", X"F3D661", X"F4D159", X"F9D45D", X"FCD462", X"FBD263", X"F8D461", X"F2D669", X"FAE588", X"A69249", X"897547", X"897853", X"7C7349", X"9B9152", X"EED776", X"EBCC5B", X"F8D163", X"FAD15F", X"F4D454", X"F4D753", X"F0D153", X"F7D772", X"E2C888", X"493612", X"201600", X"A3926C", X"FFDC8B", X"F6D162", X"EFD85B", X"F0D759", X"FCD061", X"FFC86A", X"DA8335", X"CB5E21", X"D85A2A", X"DB5B32", X"D16137", X"D05F3A", X"D65A3B", X"D05A40", X"C6684D", X"7E4332", X"291925", X"444963"),
        (X"524E62", X"1B1510", X"847342", X"F9DD89", X"F6D467", X"F9D45F", X"F8D269", X"F9D16B", X"FFD368", X"DE9744", X"BE522E", X"CF5540", X"C95632", X"BE5220", X"BA561D", X"B05011", X"BF5B16", X"C15A16", X"C4571C", X"B75A2E", X"9B5F4C", X"43201A", X"210F0A", X"A39772", X"F1DC7B", X"EAD357", X"EAD963", X"F1DA69", X"F6D160", X"FFC666", X"CF7334", X"C55530", X"CE5C43", X"C35B3A", X"CD7C3E", X"FFCB77", X"F9CF64", X"F2D35E", X"EFD55E", X"EED564", X"F6DE7B", X"BBA566", X"26170F", X"3B2B1E", X"E3CC7B", X"F4D862", X"F6D25C", X"F9D45F", X"FCD462", X"FBD261", X"F8D45F", X"F5D563", X"F6DA6D", X"F1D875", X"F4DA88", X"FDEA9A", X"E8DB86", X"F6E587", X"EBCE5D", X"F7D25A", X"FCD15D", X"FCD15D", X"F5D559", X"F4D657", X"F0D258", X"F6D975", X"E4C98E", X"493614", X"201502", X"A1926E", X"FFDC8D", X"F6D164", X"F2D65D", X"F4D55D", X"FCD061", X"FFC96A", X"D18030", X"BF5C19", X"C95922", X"CD5A2A", X"BB4E23", X"C2552C", X"CF5C36", X"D16543", X"C87254", X"743B2E", X"20081C", X"443E60"),
        (X"504F62", X"1B1510", X"847342", X"F9DD89", X"F6D467", X"F9D45F", X"F8D269", X"F8D26B", X"FFD46C", X"D69A4A", X"AE5936", X"BF5C44", X"D47543", X"D07635", X"C6742E", X"D27C32", X"D67529", X"DB7329", X"DC712F", X"D07441", X"A76D53", X"4E3122", X"211607", X"AAA478", X"F1DC7D", X"EAD359", X"ECD861", X"F2DA67", X"F4D262", X"FDC76E", X"C57447", X"B45A44", X"B05C4B", X"A45B3F", X"B67842", X"F7C574", X"F7CF68", X"F4D260", X"F2D35E", X"F1D362", X"F4DB79", X"BBA566", X"26170F", X"3D2D1E", X"E1C978", X"F4D764", X"F6D25C", X"F8D25D", X"F9D361", X"FBD462", X"F9D45F", X"F8D45F", X"F7D35F", X"F5D361", X"E3C355", X"E8CC5F", X"EBD465", X"E8CF5D", X"F6D05B", X"FBCC58", X"FCCD5B", X"FCD15D", X"F5D45D", X"F2D65D", X"EED25C", X"F2D775", X"E3CA8E", X"473514", X"1D1403", X"9E926F", X"FCDB8D", X"F4CF65", X"F4D461", X"F5D45F", X"FCD063", X"FFCB68", X"D58D36", X"C06C20", X"C86B26", X"CD6A29", X"D07234", X"CA6D36", X"C36736", X"B6643D", X"98573F", X"7E544D", X"4B3B49", X"64607A"),
        (X"504F62", X"1B1510", X"847342", X"F9DD89", X"F6D467", X"F9D45F", X"F8D269", X"F5D371", X"FFE386", X"9A7834", X"3E0C00", X"7E4528", X"FFCA85", X"FFCD6F", X"FFD068", X"FFD064", X"FFCD5F", X"FFCA61", X"FFC566", X"FFC678", X"E6C18B", X"46350F", X"211E00", X"ABA26C", X"F8DA80", X"F5CE5E", X"F5D661", X"F7DA64", X"F2D468", X"F4CC81", X"733B27", X"450D14", X"3A1818", X"381D0D", X"5D4015", X"FCDC97", X"F4D172", X"F7D263", X"F8D25D", X"F5D361", X"F5DA75", X"B9A462", X"271910", X"3F2F20", X"DFC877", X"F5D865", X"F7D35F", X"F7D15C", X"F7D15C", X"FED863", X"FFD966", X"FAD15F", X"FAD05C", X"FDD05B", X"FFD55B", X"FFD659", X"F9D557", X"F6CF56", X"FFD064", X"FFCC63", X"FFCB5E", X"FDD05F", X"F4D461", X"F0D661", X"EDD35C", X"EFD774", X"E2CC91", X"453616", X"1B1503", X"9D9271", X"FADC8F", X"F4CF67", X"F6D162", X"F7D060", X"FCD063", X"FFCD66", X"FFCB6B", X"FFC86D", X"FFC770", X"FFC770", X"FFC96C", X"FFC877", X"FFC78D", X"6D3E1E", X"290801", X"9F8F92", X"FFFFFF", X"F2FDFF"),
        (X"504F62", X"1B1510", X"847342", X"F9DD89", X"F6D467", X"F9D45F", X"F8D269", X"F3D371", X"FAE58A", X"917B3A", X"2E1200", X"6E4C2C", X"F9D181", X"FDD467", X"F7D662", X"F7D75E", X"F9D559", X"FED25B", X"FFCC5F", X"FDCC72", X"DEC687", X"413809", X"1E2100", X"AAA368", X"F8DA7C", X"F6CD5E", X"F6D561", X"F8D966", X"F3D768", X"EECE7B", X"68401E", X"401D12", X"352216", X"2F2106", X"604614", X"F4D289", X"F7CF72", X"FAD063", X"FAD25D", X"F7D261", X"F3D972", X"B9A462", X"27190E", X"403021", X"DEC776", X"F7DA66", X"F8D461", X"F6D05B", X"F1CE56", X"FFDF69", X"FFE073", X"FCCD64", X"FDCA60", X"FFD061", X"FFD059", X"FFCA4D", X"FCCA4E", X"FFCD5A", X"FFBF65", X"FFC06A", X"FFC763", X"FFCE61", X"F4D461", X"EFD761", X"EDD35C", X"EED671", X"E2CE90", X"423613", X"191500", X"9C916E", X"F8DC8C", X"F3CD66", X"F7D062", X"F9D060", X"FCD061", X"FDCF61", X"FFCE65", X"FFCE65", X"FFCE66", X"FFCE66", X"FFCF62", X"FBD06D", X"F0CF8D", X"5B4622", X"190E0D", X"94929E", X"FBFFFF", X"F2FEFA"),
        (X"505060", X"1B1510", X"847342", X"F9DD89", X"F6D467", X"F9D45F", X"F8D367", X"F3D46F", X"FCE584", X"917D34", X"271500", X"674F2E", X"F7D27F", X"FCD469", X"F7D568", X"F6D666", X"F6D55F", X"F9D45F", X"FFCD63", X"FACD78", X"DCC68B", X"3E390D", X"1B2100", X"A5A668", X"F1E074", X"EDD456", X"F3D665", X"F7D96A", X"F2D561", X"E9CE61", X"DBBC63", X"CBAB64", X"D1B278", X"D3B073", X"D8A95E", X"FFD179", X"FFCC66", X"FFCE5F", X"FCD05F", X"F5D266", X"F3D874", X"B9A560", X"281A0F", X"413122", X"DEC776", X"F8DB67", X"F9D562", X"F6D05B", X"F3D154", X"FDD961", X"E6BC54", X"B98628", X"BD8027", X"F3AF54", X"FFC863", X"FFC75C", X"FFC45A", X"FABA5E", X"C87C3D", X"BE7135", X"FFC56B", X"FFCE61", X"F5D361", X"EFD75F", X"ECD55B", X"EDD76F", X"E3D090", X"42360F", X"191600", X"9A936A", X"F8DC8A", X"F3CE62", X"FACF60", X"FCCF5C", X"FCD15D", X"FCD15D", X"FDD25D", X"FDD25D", X"FCD45E", X"FED45E", X"FFD25E", X"F9D16B", X"EBD387", X"554A1E", X"15110D", X"9292A2", X"FFFFFF", X"FAFAFE"),
        (X"524F60", X"1D140E", X"85733E", X"F9DE85", X"F6D463", X"F9D45D", X"F8D365", X"F5D36F", X"FDE388", X"8F7D38", X"241600", X"664F32", X"FACF87", X"FFD06F", X"FCD16E", X"F9D46A", X"F6D463", X"F9D363", X"FFCC68", X"FACC7A", X"DCC68D", X"3E3911", X"1B2100", X"A3A66C", X"F1DF78", X"EDD35A", X"F2D56B", X"F5D96E", X"EED65C", X"EBD556", X"F2DA63", X"FDE178", X"FFE08C", X"FFD785", X"FFD578", X"FFD169", X"FFCC5C", X"FFCE5D", X"FCD063", X"F5D26A", X"F3D874", X"B9A560", X"271B0F", X"403222", X"DEC776", X"F9DA69", X"F7D664", X"F4D15B", X"EFCA4E", X"FFD966", X"F6BC60", X"BD782B", X"B76624", X"FFAE69", X"FFD181", X"FFC670", X"FFBC68", X"FFB36E", X"C4653A", X"BF6536", X"F1B159", X"FDD163", X"F5D45F", X"F0D65D", X"ECD55B", X"EDD76F", X"E1D18E", X"42370D", X"191600", X"9A9466", X"F6DE84", X"F3CF60", X"F9D05E", X"FAD05C", X"FCD05F", X"FDD05F", X"FFD061", X"FFD063", X"FFD064", X"FFCF66", X"FFCC68", X"FFCC75", X"EED08F", X"574824", X"151011", X"9491A4", X"FFFDFF", X"FEF7FF"),
        (X"554D60", X"20130C", X"87733A", X"FADF7F", X"F6D65D", X"FBD457", X"FBD263", X"F8D073", X"FFE394", X"8C7642", X"1A0A00", X"583A2B", X"D89B69", X"DF994F", X"FFCF7B", X"FFD371", X"FAD161", X"FCD061", X"FFCC68", X"FCCB7A", X"DEC58D", X"413711", X"1E1F00", X"A8A270", X"F8D886", X"F5CC68", X"F3D371", X"F2DA6E", X"E7D555", X"E8D953", X"F5E068", X"E7C95D", X"F1C267", X"FAC76B", X"F8CA61", X"F3CA58", X"F8CF5B", X"FAD15F", X"FAD066", X"F7D16C", X"F5D776", X"B8A560", X"241D0F", X"3C3422", X"E0C678", X"FBD969", X"F6D664", X"F4D15B", X"F1C751", X"FFCF68", X"FFB56A", X"C05B27", X"CD5E34", X"E7724A", X"F48954", X"ED854A", X"F78F57", X"F18354", X"D25538", X"C55D30", X"F0BB5D", X"F3D75F", X"F9D85F", X"F5D65D", X"EFD55C", X"EED870", X"E2D28F", X"43380E", X"1A1800", X"9B9565", X"F7E07F", X"F3D25B", X"F5D45F", X"F7D261", X"FCCF66", X"FFCB6A", X"E7A54E", X"D18538", X"DA8641", X"E38A48", X"E38A48", X"DB8E56", X"CE9876", X"5D3A2F", X"291822", X"A196AC", X"FFF9FF", X"F1E9FE"),
        (X"534E60", X"1E140C", X"87733A", X"FADF7F", X"F6D65D", X"F9D557", X"F9D363", X"F5D371", X"F8DC8C", X"826D37", X"1B0D00", X"52351F", X"9F602F", X"AC611B", X"F9BC66", X"F7C561", X"FAD15F", X"FAD15F", X"FFCC66", X"FCCC78", X"DEC58B", X"41370F", X"1E1F00", X"A8A270", X"FAD788", X"F6CB6A", X"F5D36F", X"F3DA6A", X"E4D04C", X"F2DD57", X"FFE570", X"FFDC74", X"FFD278", X"FFD77C", X"FFD56B", X"EDCA56", X"F5D45D", X"F7D35F", X"FAD066", X"F8D06C", X"F3D876", X"B5A760", X"1F1F0F", X"383622", X"DEC778", X"F9DA69", X"F4D764", X"F1D25D", X"F8CF5D", X"FFCC69", X"FFB774", X"CB6C3F", X"BF4F33", X"CC553D", X"C75230", X"CC5733", X"C7522E", X"D25C3D", X"C54C35", X"C16235", X"EBBD5D", X"F3D960", X"FDD760", X"F9D45D", X"F1D55C", X"EED872", X"E4D191", X"43380E", X"1A1800", X"9B9663", X"F9E07D", X"F3D259", X"F2D65B", X"F4D45F", X"F8D166", X"FFCC6C", X"C17C28", X"AF5D17", X"B4581A", X"B3541B", X"B5551E", X"AA5627", X"9D6040", X"441B0B", X"1B0201", X"998995", X"FFF8FF", X"FFF6FF"),
        (X"4B525E", X"18170E", X"84733E", X"F9DE85", X"F5D563", X"F6D65B", X"F3D663", X"F0D66D", X"F2DF7F", X"9E8F42", X"584F1B", X"745F2D", X"B7853D", X"C38930", X"FBCC65", X"FCD565", X"F5D45B", X"F7D45B", X"FFCE61", X"F8CE74", X"DBC887", X"3E3A0B", X"1B2200", X"A5A56A", X"F5DB80", X"F3CE62", X"F3D567", X"F7DA64", X"EFD14C", X"FCD654", X"EFBB4D", X"EEB053", X"F2AF60", X"EBAE5C", X"ECBA59", X"F6CD60", X"F8D25F", X"F8D261", X"FCCF68", X"F8D06C", X"F0DA74", X"B0AA5E", X"1A210F", X"333922", X"DAC978", X"F6DB69", X"EFDA64", X"EBD55F", X"F3D665", X"FCD875", X"E6BC73", X"955E2C", X"9B4E31", X"BE5D4C", X"CD5745", X"CC4D3C", X"CF5442", X"C95A49", X"9E4833", X"925326", X"E6BF61", X"F9D763", X"FFD460", X"FFD15D", X"F4D25E", X"EFD676", X"E6D093", X"453710", X"1B1700", X"9D9465", X"FADF7F", X"F3D259", X"EFD857", X"EFD859", X"F4D55D", X"FAD161", X"D19B37", X"C9882F", X"D38836", X"CE7F35", X"C87D39", X"BD7A3A", X"B38243", X"845F2C", X"5F4424", X"9B867A", X"D5BFCB", X"DAC2DA"),
        (X"48545E", X"14150C", X"857144", X"FCDB8F", X"F8D26D", X"F8D461", X"F2D665", X"EDD869", X"ECD970", X"E4D477", X"E3D68D", X"FCE69E", X"FBD076", X"FFD068", X"F9D060", X"F7D35D", X"F5D559", X"F8D35B", X"FFCE61", X"FACD74", X"DCC689", X"3E3A0B", X"1F2600", X"A6A568", X"F5DC7A", X"F3CF5C", X"F6D465", X"FBD864", X"FED556", X"FDC74E", X"C17B18", X"AD5C0C", X"B66324", X"A55616", X"C0832D", X"FCCB67", X"FAD063", X"F8D163", X"FAD068", X"F5D16C", X"F0DA74", X"B0AA5E", X"1A210F", X"303620", X"DAC978", X"F6DB6B", X"EFD966", X"EBD561", X"EBD262", X"FDE685", X"CAB96F", X"4A3000", X"481700", X"974941", X"C75857", X"CB5050", X"CC5758", X"A64944", X"521B0C", X"330F00", X"E2C069", X"FDD668", X"FFD262", X"FFCF5F", X"F7D062", X"F3D478", X"E7CE97", X"483414", X"1F1500", X"A09267", X"FCDD83", X"F4D15B", X"F0D759", X"EFD857", X"F2D65B", X"F7D35D", X"FCCE60", X"FFC963", X"FFD676", X"FFCE77", X"FFD081", X"FFCB7E", X"FDD07D", X"E9C578", X"FDDFA7", X"947B5D", X"1A0004", X"52384C"),
        (X"4A535E", X"171310", X"836645", X"FDD094", X"FCC873", X"FACB64", X"F0D165", X"EFD86A", X"F3DA6C", X"F2D871", X"E9D275", X"F0D276", X"FACF6A", X"FDCF61", X"F6CE5C", X"F6D05B", X"FBD35F", X"FFD869", X"FFD06B", X"F7C272", X"DBBD88", X"493A14", X"292603", X"ADA46E", X"FFDE7E", X"FED161", X"FFD669", X"FFD96B", X"FFD662", X"FFC95C", X"CC7C2A", X"BA5C1E", X"CE6239", X"C15B2E", X"C97935", X"FFC870", X"FCCF68", X"F5D363", X"F4D366", X"F0D46A", X"F8E37A", X"B9AC63", X"1C1F0C", X"353420", X"DAC273", X"F5D467", X"F0D261", X"E9CE5F", X"EBCE64", X"F3DE81", X"C9C27E", X"372E04", X"3B210E", X"894F51", X"C26270", X"BC5062", X"B75967", X"904D54", X"3A1F18", X"3E2F0D", X"D3B468", X"FFD671", X"FFCB62", X"FFCB60", X"FACE66", X"EFCB75", X"E7C897", X"4D331A", X"261705", X"A5926E", X"FED986", X"F5CC5D", X"F7D861", X"F5D961", X"F9D861", X"FCD663", X"F6CB5A", X"FDCA5E", X"FFC961", X"FFC665", X"FDC56F", X"FECA72", X"F5C767", X"EFC76B", X"F9DA92", X"8D7448", X"26100A", X"5A4855"),
        (X"575C68", X"201516", X"6C422B", X"B57649", X"C57F39", X"FFC26A", X"F7CF68", X"EFCE63", X"FBD66A", X"FCD26A", X"F5CD66", X"FACF6A", X"FDCF63", X"FFCE61", X"FACC5E", X"FCCC61", X"FFCB64", X"FFD172", X"F6AD58", X"BA7534", X"AB7D55", X"442811", X"2E1C09", X"B59C72", X"FFCF79", X"FDC359", X"FEC866", X"FFCC6A", X"FFCF67", X"FFC164", X"C77533", X"B65428", X"C95C3F", X"BE5433", X"C67336", X"FFC171", X"FFCE6B", X"FBD167", X"FBD167", X"F8D269", X"F7D571", X"BBA55C", X"261D0E", X"403525", X"E5C378", X"FFD56D", X"FBD368", X"F4CF65", X"E4BE59", X"FCDE8B", X"D2C78D", X"302A07", X"321F18", X"491E2A", X"63162E", X"63112C", X"58192F", X"4D2633", X"2C2225", X"342F15", X"D0B470", X"FFD677", X"FFCB66", X"FFCC64", X"F3C663", X"FBD282", X"EFCAA0", X"4F331F", X"29170B", X"A58C6E", X"FFD78A", X"FFCE69", X"FCD268", X"FBD368", X"FCD268", X"FED266", X"FAC95F", X"FFCC62", X"FFCC63", X"FFC764", X"FEC76C", X"FFCA70", X"FAC664", X"F3C76B", X"FBDA8E", X"8F7749", X"24190D", X"595458"),
        (X"554E5C", X"260E14", X"71352C", X"B05D3E", X"CB7038", X"FFC174", X"FFD373", X"FFE079", X"FFD672", X"FFD170", X"FFCC68", X"FFD069", X"FFD06B", X"FFD06D", X"FFCC6C", X"FFCC6F", X"FFCC77", X"FFCC81", X"FFA362", X"BE6639", X"A2614E", X"512220", X"320D0E", X"C1957F", X"FFCA85", X"FFBE65", X"FFC672", X"FFCB79", X"FFD67E", X"FFCA7D", X"CA7E4D", X"B55F41", X"C56954", X"BB6243", X"C97E45", X"FFC97E", X"FFCF73", X"FFCF6B", X"FFCD6B", X"FFCD6D", X"FFD575", X"CAA260", X"311A0F", X"4B3025", X"F2C27C", X"FFD471", X"FFD26B", X"FFCE69", X"FFD378", X"FFE097", X"DCBF90", X"3F2915", X"361F24", X"351128", X"3E0725", X"3E0C2A", X"341B33", X"2B2135", X"35303D", X"302619", X"D8BE80", X"FFE187", X"FFD875", X"FFD773", X"FFD373", X"FFD990", X"EAC09A", X"573525", X"270E09", X"AE9279", X"FFDD94", X"FFCB6C", X"FFD57A", X"FFD47C", X"FFD57A", X"FFD377", X"FFD275", X"FFD474", X"FFD573", X"FFD273", X"FFD077", X"FFD47C", X"FFCF75", X"FFD07D", X"FFDB9A", X"88764A", X"111501", X"404D46"),
        (X"665F6D", X"2E131C", X"793736", X"C36857", X"C35D32", X"DA7A38", X"D28838", X"D5913D", X"DB8A3D", X"DE8639", X"D9802F", X"DB8432", X"D88536", X"D68638", X"D58137", X"D9803C", X"E6844A", X"E7804C", X"D56B3A", X"B35432", X"9E5950", X"4B181B", X"380B14", X"AB7265", X"E28751", X"E07A32", X"DE803E", X"DC8646", X"E39854", X"D38F57", X"874A2C", X"6A2F1F", X"773B2F", X"71321E", X"8C471F", X"D98E56", X"D4823C", X"D98232", X"DE802C", X"D98230", X"D18C3D", X"A06D3A", X"2A100B", X"4B2927", X"C27D4B", X"E08D42", X"DB8B3B", X"D58738", X"DA8A45", X"D18D56", X"B68968", X"402419", X"392530", X"4A344E", X"614062", X"614568", X"38314F", X"22253D", X"343346", X"30211D", X"A2774A", X"D29951", X"CD923D", X"D0903B", X"D48E44", X"D6915B", X"C0876D", X"52241B", X"371613", X"88604E", X"CA8B51", X"D08337", X"D5853E", X"D68440", X"D6853E", X"D6853C", X"D6853A", X"DA893C", X"DA8C3B", X"D98839", X"DC863B", X"DF8A40", X"DA833C", X"D18445", X"D29C6C", X"674A2B", X"19180D", X"3B4949"),
        (X"494F58", X"190913", X"69303A", X"BF6964", X"CD6542", X"C95B27", X"C05925", X"BD5323", X"C65227", X"CB5027", X"CB5025", X"CB5025", X"C95027", X"C95027", X"C64D24", X"C74B2A", X"CD4A36", X"CE503B", X"CB5A37", X"C46A4B", X"A0675D", X"492020", X"371012", X"7F4136", X"C2542E", X"D24F1E", X"CF5022", X"CA5226", X"C5582B", X"AB5A38", X"4C251A", X"251516", X"2E1E1F", X"391A17", X"66261C", X"B95C47", X"C25430", X"CA5320", X"C95616", X"C1591A", X"BC6636", X"874E34", X"2B181E", X"472732", X"B25245", X"C84C2D", X"C54E29", X"C44F29", X"C8502F", X"B8533A", X"8F5444", X"40231D", X"352D34", X"312D43", X"3C2D50", X"3F3057", X"262145", X"232341", X"222539", X"351E21", X"A65A48", X"BA552E", X"BA581E", X"BD561E", X"C6512D", X"C1503D", X"AB534A", X"5F1D1D", X"471518", X"864A43", X"BD603D", X"C25322", X"C24F22", X"C44E22", X"C24F22", X"C04F1E", X"BF4E1B", X"BF521C", X"BF541B", X"BE511A", X"C14E1E", X"C65024", X"C24A1E", X"B94B25", X"AB563E", X"6B342B", X"25131E", X"525166"),
        (X"788388", X"68626B", X"865D6D", X"8B454D", X"9C3D29", X"C95B39", X"D25C3B", X"CB4E2F", X"D9543B", X"DA533D", X"DA533D", X"DA533D", X"DA533D", X"DA533D", X"D75039", X"DA4F3E", X"E3524E", X"D44E49", X"B64F39", X"893F2A", X"794949", X"3B1721", X"351016", X"955751", X"CE5C45", X"E25537", X"E05539", X"DB573B", X"D65D41", X"B9614F", X"513034", X"232330", X"202533", X"2C1F28", X"63272B", X"BB5C56", X"CB513F", X"D34F31", X"D15227", X"C8562D", X"C06048", X"894A42", X"2B1724", X"482837", X"C0575B", X"D84F44", X"D5523E", X"D3533E", X"D75347", X"C65850", X"9D5A53", X"472727", X"251D27", X"29283D", X"33294C", X"2D224A", X"252147", X"232343", X"222539", X"3A1D26", X"BB5D5D", X"D15647", X"D15937", X"D45835", X"D34B3A", X"CD4E47", X"B25250", X"661F22", X"430C13", X"894747", X"CB644E", X"D8593B", X"D95539", X"DA5437", X"D95537", X"D65533", X"D35530", X"D45930", X"D45B32", X"D15831", X"D65437", X"DD563D", X"D95035", X"CE523A", X"BF5F52", X"78383A", X"270F23", X"4C4764"),
        (X"F2FDFF", X"F9FAFF", X"A892A9", X"24000C", X"6E2529", X"B9594E", X"CA5541", X"CC4E34", X"D4573D", X"D2573F", X"D2573F", X"D2573F", X"D2573F", X"D2573F", X"CF533B", X"D3533E", X"E3594F", X"CD554E", X"9A5040", X"3C0A04", X"441931", X"391131", X"3C1929", X"864D50", X"C65D55", X"D65749", X"D55849", X"D25949", X"D15D4B", X"B95F59", X"552C3C", X"291E38", X"20233B", X"29202E", X"5C2A2D", X"B55F58", X"C55441", X"CE5137", X"CE5135", X"C8533D", X"BF5F54", X"8C4848", X"311422", X"4E2535", X"BB5A59", X"CF5346", X"CB573E", X"CA573E", X"CE574B", X"C15956", X"9D5957", X"4C2529", X"36212F", X"64556C", X"6D5579", X"3C284C", X"252241", X"22243F", X"252439", X"3B1B2A", X"B95C65", X"CF5553", X"D25645", X"D4563F", X"CF4E38", X"C55343", X"A8584E", X"5E2224", X"3B0E19", X"84484D", X"CA6354", X"D65841", X"D7543F", X"D7553D", X"D6563D", X"D35639", X"D05636", X"D15937", X"D05B38", X"D05739", X"D45343", X"DB5547", X"D4513B", X"C7553E", X"BE6858", X"77403E", X"281529", X"4E4E6C"),
        (X"F0FEF9", X"FAFFFF", X"ADA8B7", X"422A3D", X"5A2A38", X"9C595D", X"A14C42", X"B35444", X"B35547", X"B35547", X"B35547", X"B35547", X"B35547", X"B35547", X"AF5244", X"B25247", X"B5524A", X"AD5C55", X"7A4B44", X"2F0E12", X"421A33", X"3E1737", X"2F1229", X"774E5C", X"A7595F", X"B25555", X"AF5755", X"AF5753", X"B25A51", X"9E5A5C", X"43233E", X"1A1436", X"1E233C", X"262132", X"502D32", X"A2635F", X"AE5851", X"B6554B", X"B6554D", X"B15653", X"AF6366", X"814B54", X"2E1428", X"482739", X"9F575D", X"AC544D", X"A95747", X"A95747", X"AE5650", X"A55758", X"875558", X"3C1D26", X"271426", X"352640", X"3D2848", X"2C1D3D", X"23233F", X"1E263F", X"22253D", X"331E33", X"9B5969", X"AD535A", X"B05350", X"B2544A", X"B15647", X"A9594D", X"965B58", X"4E2429", X"391928", X"784D57", X"AE625A", X"B35444", X"B44F46", X"B44F46", X"B35046", X"B05043", X"AD5040", X"AE5440", X"AD5641", X"AE5143", X"B34D4B", X"B84F4E", X"B14C42", X"A64F41", X"A6665C", X"6A4443", X"2C202D", X"5C5E72"),
        (X"EEFFF7", X"E8FAED", X"F0F5F1", X"FFFFFF", X"C9B7C2", X"351D27", X"3D2325", X"4A292B", X"472026", X"491E28", X"491E28", X"491E28", X"491E28", X"491E28", X"451B25", X"421D23", X"3D2222", X"3B2624", X"3A292D", X"41292F", X"8E6469", X"512834", X"36243E", X"3B2B49", X"4D2B42", X"44202E", X"41222A", X"422425", X"441D1D", X"4A2D37", X"201D3E", X"2D375C", X"1B243C", X"212332", X"2F1F2B", X"381B25", X"441B27", X"491E2A", X"461D2D", X"452031", X"422231", X"392434", X"2C2840", X"2D263F", X"3A2032", X"43212C", X"3F2328", X"412326", X"432025", X"402127", X"35262D", X"2C2734", X"26273B", X"252842", X"272541", X"22223F", X"1E2541", X"1E2943", X"1C2A45", X"242641", X"342135", X"391E2C", X"391F28", X"432C2F", X"392125", X"3B2329", X"3F262F", X"342030", X"352841", X"38273B", X"432627", X"492221", X"4A2029", X"4B1D2C", X"491E2A", X"461E27", X"431E24", X"442126", X"442327", X"442126", X"421924", X"522431", X"52232E", X"481E25", X"3B1D20", X"9D8A8E", X"FFFFFF", X"F1F2F6"),
        (X"F4FFF6", X"EDFDEF", X"F0FBF1", X"EEF3F1", X"D5D5DE", X"27232B", X"201D17", X"261F13", X"2D1E16", X"2F1E16", X"2F1E16", X"2F1E16", X"2F1E16", X"2F1E16", X"2B1A12", X"291D11", X"21210A", X"25240C", X"2F2212", X"422B23", X"9C7876", X"4E2E39", X"251C38", X"20203B", X"1B121E", X"2F2625", X"29291D", X"2A2816", X"31220C", X"24160A", X"1F212E", X"364058", X"1C2737", X"1F2633", X"252233", X"282133", X"332738", X"302232", X"221822", X"281F22", X"2B1E1A", X"2A2018", X"252120", X"221F25", X"282027", X"2C242E", X"28242E", X"262123", X"261F11", X"251D09", X"221E0D", X"1E1D12", X"1C1B17", X"1E1C1A", X"1E1A19", X"191713", X"151B14", X"141E19", X"131E1F", X"141D1F", X"252623", X"292822", X"2A2923", X"161712", X"292F33", X"1F2125", X"2B201D", X"1F120B", X"24201D", X"24201B", X"2A1F0E", X"2C1C0D", X"2E1A15", X"2E1816", X"2D1916", X"2A1913", X"271910", X"281C10", X"271E11", X"261D12", X"261C14", X"271C1B", X"2F2029", X"3A2C3A", X"180D1A", X"9B959B", X"FAFDF5", X"EFF6E8"),
        (X"FFFEF9", X"F9FAF7", X"F6FFFF", X"CCD6DC", X"4D5160", X"2D282A", X"9A8B69", X"B29F68", X"B4A364", X"B4A360", X"B4A360", X"B4A360", X"B4A360", X"B4A360", X"B0A05D", X"B3A15C", X"B4A055", X"BAA256", X"C1A15C", X"A8885E", X"462E32", X"3A2C45", X"34374F", X"151921", X"716953", X"B1A87B", X"A7A971", X"A5A463", X"B3A15A", X"BCA468", X"BAA988", X"615A4F", X"1F2827", X"1C2733", X"1F243B", X"222339", X"2A2836", X"2A2622", X"878568", X"B9B483", X"B7A269", X"BBA165", X"BAA06D", X"B7A077", X"AD9C84", X"4B3F33", X"241B17", X"6A624E", X"B1A96C", X"B4AA5C", X"B7A860", X"B8A562", X"BAA165", X"BDA169", X"BDA065", X"B3A060", X"ABA65F", X"A8AA65", X"ABA76D", X"ADA671", X"ACA36D", X"B3A772", X"BAA978", X"796A49", X"241C11", X"453E31", X"B1A479", X"AEA264", X"ACA465", X"AEA463", X"B4A163", X"B89D62", X"B99C64", X"BA9A63", X"B89B63", X"B69B5F", X"B39B5C", X"B49E5D", X"B3A05E", X"AFA05F", X"ADA867", X"989566", X"383327", X"221F27", X"7B7B8B", X"D4D7DF", X"F8FFF1", X"EFFADD"),
        (X"FFFBFF", X"FFFBFF", X"FDFFFF", X"BAC1C1", X"0A0701", X"31230A", X"DDC383", X"FFE892", X"FEE283", X"FCE381", X"F9E57F", X"F8E67F", X"F8E67F", X"F9E57F", X"F7E17B", X"FCE17A", X"FEDF73", X"FFE077", X"FFE07D", X"EFC881", X"271100", X"19141A", X"1F2430", X"0E110B", X"95885D", X"F6E6A0", X"EAE68F", X"E6DF7D", X"EBD771", X"F3DB7F", X"FCE6A7", X"706341", X"222821", X"1C2733", X"1D253D", X"1F243D", X"252C39", X"1F2317", X"B7B781", X"EEE594", X"F3DA81", X"F9D87B", X"FBD681", X"F6D68F", X"ECDCA8", X"5D5233", X"1C1007", X"887A5F", X"F5E592", X"FCE77A", X"FFE57C", X"FFE17F", X"FFDE80", X"FFDD83", X"FFDC82", X"FEDB7C", X"F4E379", X"F3E77E", X"F6E386", X"F8E18C", X"F0D984", X"F8E18E", X"FEE69A", X"9B8954", X"1B1202", X"4E4632", X"EEDE9A", X"F5E284", X"F0E27E", X"F3E17E", X"F9DD80", X"FDD981", X"FDD981", X"FCD880", X"FAD97E", X"F7D97B", X"F6D877", X"F7DC7A", X"F6DE79", X"F2DE7A", X"F3E785", X"DCD585", X"3D360D", X"181609", X"BDC0C8", X"F1FBFF", X"FCFFF8", X"FAFFEC"),
        (X"FFFDFF", X"C7C8D0", X"939894", X"8E8B75", X"7C6637", X"A17F39", X"E7C264", X"FBD36A", X"F3C75F", X"F8D068", X"F3D866", X"EBD55F", X"EAD760", X"E0C752", X"F5D363", X"F7D060", X"F7D15C", X"F9D05C", X"FACE62", X"F6CE70", X"8D7229", X"7D7042", X"38382D", X"0D0800", X"A08654", X"FDDF8E", X"E5CE69", X"E9D764", X"EAD963", X"E1D26A", X"ECDD90", X"6D6437", X"0E140D", X"333949", X"2E2F45", X"22253D", X"1F2B40", X"162016", X"AAA462", X"F9E686", X"EED36A", X"F2D266", X"F2D266", X"ECD372", X"E0D58E", X"564D22", X"1A0C01", X"907B65", X"FFDC8D", X"F8D163", X"F2CE5D", X"F8D463", X"FDD66A", X"F6CC64", X"FBCB6B", X"FFD471", X"F3CE62", X"F0D060", X"F0CF64", X"F2CE68", X"F2CC67", X"E7C865", X"F5E189", X"8D8346", X"121003", X"453F2F", X"E7D187", X"EFD368", X"F0D769", X"F2D667", X"F8D367", X"F9D267", X"F4CF67", X"EFCC64", X"E9C65E", X"EECD62", X"EFCF61", X"EBCE5D", X"EBCE5D", X"ECD15F", X"F3DB68", X"E8D26C", X"8C7929", X"726837", X"898D85", X"98A5AA", X"B6C2BE", X"F6FFFA"),
        (X"F9FDFF", X"6D6F7A", X"080B05", X"605738", X"FFEBA6", X"FFE182", X"FFD667", X"F6C956", X"FFCE61", X"FBCB5E", X"F8CF5F", X"FCD663", X"FFDA68", X"FFD866", X"FFD568", X"FECE5E", X"F9CF57", X"FAD058", X"FCCE5E", X"F7D064", X"FEE17E", X"ECDC94", X"54513B", X"251C0D", X"A58452", X"FFDB8A", X"EDCC61", X"EFD55C", X"ECD95D", X"E1D364", X"ECDE88", X"6D6631", X"0C0C08", X"3D3E52", X"38344C", X"1C1D36", X"1E2945", X"171E1C", X"AEA35E", X"FDE67C", X"F1D362", X"F2D35E", X"F4D25E", X"EFD26C", X"E4D588", X"574D1E", X"1B0D02", X"927A65", X"FFDB8D", X"FAD161", X"F4CE57", X"F9D45D", X"FBD35F", X"FFCE63", X"FFCC6B", X"FFCA6D", X"FFCC69", X"FFCD69", X"FFCE6C", X"FFCE6C", X"FFD776", X"FFCF72", X"FADD89", X"978953", X"13100A", X"464032", X"EAD284", X"F2D362", X"F5D563", X"F6D561", X"FBD35F", X"FDD261", X"F2C85D", X"FFDE77", X"FCCD66", X"FFD36B", X"FFD166", X"FDD465", X"F4D260", X"EECF5A", X"F2D15A", X"F4D463", X"F7DC7A", X"F7E7A4", X"5A5C4C", X"000207", X"727D80", X"F6FFFF"),
        (X"F8FCFF", X"777A84", X"101211", X"5D5438", X"F1D18A", X"F5CA67", X"F8CD5E", X"F9CE5B", X"FBCD5F", X"FFCD63", X"FFC866", X"FFBF63", X"FFB85F", X"FFBA60", X"F4B657", X"FBC55F", X"FCCF5A", X"FAD058", X"FCCE5E", X"F7D064", X"EED16D", X"E7D78F", X"423F2A", X"20170A", X"A88256", X"FFD98E", X"F0CA63", X"F2D45C", X"EFD75D", X"E4D262", X"EFDE84", X"72632F", X"160F0F", X"3A3650", X"322E46", X"24213D", X"222649", X"1C1B20", X"B2A160", X"FFE57C", X"F1D460", X"F4D35C", X"F9D060", X"F6CE70", X"ECD08C", X"5C4A20", X"1D0D00", X"907C61", X"FBE08C", X"F3D663", X"EED358", X"F7D75E", X"FBCE5B", X"FFCF67", X"FFC76B", X"FFB865", X"FFB364", X"FFB369", X"FEB36B", X"FFB26B", X"FFBD76", X"FEB774", X"F2BE85", X"A28360", X"1A1112", X"4A4335", X"EDD687", X"F6D666", X"F5D563", X"F6D561", X"FBD35F", X"FED063", X"FCCA69", X"FDC069", X"FAB25D", X"FFB45E", X"F9B158", X"FFC86A", X"FFD872", X"F1D163", X"FAD663", X"EDCB5B", X"EACA69", X"EDDB98", X"626353", X"0F171D", X"82888D", X"F8FEFF"),
        (X"FAFFFF", X"7C7F89", X"0A0C0E", X"5D543A", X"F3D48A", X"FFD772", X"FED264", X"FACF5E", X"FFD767", X"FFD36B", X"EDA24E", X"BD631B", X"C96925", X"BF631E", X"B1671A", X"DCA043", X"FCCE5E", X"FAD058", X"FCCE5E", X"F7D064", X"EED16D", X"DDCD85", X"4D4A34", X"23170E", X"AB7F5A", X"FFD594", X"F5C767", X"F3CF5C", X"F1D55A", X"EAD15F", X"F5DE7F", X"776327", X"2C1C19", X"30253B", X"251F35", X"34304B", X"292441", X"241918", X"B5A05C", X"FFE57A", X"F2D65D", X"F6D059", X"FFCC62", X"FEC974", X"F4CB92", X"624622", X"200C00", X"928160", X"F6E38A", X"F0D863", X"EDD358", X"F7D75E", X"FFD663", X"FDC15A", X"DE9237", X"B85D13", X"C36024", X"C55E2A", X"C35E2C", X"C35E2E", X"C85D2F", X"C15F35", X"B86C48", X"7B4A36", X"23151A", X"443D30", X"E8D081", X"F0D060", X"F5D563", X"F6D561", X"FBD35F", X"FFD063", X"EEB158", X"B3691C", X"C1671C", X"C16119", X"B35B0D", X"E39C47", X"FFD372", X"F6D56C", X"FBD462", X"FFD96C", X"EFCA6C", X"F9E1A0", X"686355", X"050810", X"76787E", X"FFFFFF"),
        (X"FDFFFF", X"7F828A", X"0E0F15", X"615741", X"FADC8D", X"F8CE63", X"FFD367", X"FBD263", X"F8D463", X"FFD771", X"F5A159", X"C05621", X"C04E23", X"C95F30", X"BC662A", X"F4B262", X"FECD60", X"FAD05A", X"FCCF5C", X"F7D064", X"F5D872", X"E0D088", X"4B4732", X"1E0F09", X"B88669", X"FFD9A1", X"F9C36B", X"F8CD5C", X"F7D459", X"EFD059", X"FCDF79", X"7A611C", X"2C1703", X"30212A", X"29233A", X"342E44", X"382A36", X"3B2610", X"B79D4F", X"FFEA78", X"F2D757", X"F9D158", X"FFD36F", X"FFBB72", X"F7C191", X"6E4729", X"271000", X"95845E", X"F8E48B", X"F1D964", X"EED559", X"F9D85F", X"FFD562", X"FFC962", X"D78B30", X"BC5C16", X"D0582C", X"D55434", X"D55336", X"D55338", X"D55137", X"CB503A", X"C85F50", X"88423E", X"29131D", X"433C2E", X"E6CF80", X"EFCF5F", X"F4D461", X"F5D45F", X"FAD25D", X"FFCD61", X"F5AC57", X"B86017", X"C6621B", X"C9621C", X"B75A0F", X"E9A04C", X"FFD473", X"F4D36A", X"FAD15F", X"FDCF63", X"F4CA6D", X"F8D99A", X"6B6054", X"0E0C16", X"7E7B83", X"FFFFFF"),
        (X"FEFFFF", X"7F828A", X"0E0E19", X"615643", X"FADC8B", X"F8CF5F", X"FFD367", X"F9D363", X"F6D762", X"FFD772", X"ED9D5D", X"B74E26", X"D05C41", X"CD5D41", X"B95D2F", X"F1A861", X"FFCC64", X"FAD05A", X"FCCF5C", X"F7D062", X"F5D872", X"E0D186", X"4B4734", X"1E0E0D", X"89513D", X"C98354", X"D69B48", X"FFD266", X"FFD75C", X"F2CF55", X"FFE175", X"CDAE60", X"C8AF88", X"94837B", X"1B162A", X"322B3B", X"AF9B8B", X"CCB37E", X"F3D77A", X"FFE66E", X"EDD04C", X"FFD659", X"FFC165", X"CD7C3C", X"C5825D", X"66351F", X"2E1603", X"907E55", X"FDE38A", X"F5D865", X"F1D55A", X"FAD960", X"FFD361", X"FFCC63", X"D69134", X"C0651D", X"D0592F", X"D85339", X"D8533B", X"D8533D", X"DC5440", X"CE4F3F", X"CD6158", X"944B4C", X"2A1420", X"453E31", X"E9D183", X"F1D161", X"F4D461", X"F5D45F", X"FAD25D", X"FFCC61", X"FDAE57", X"B85A0F", X"C35D12", X"FB9B4C", X"FFAD58", X"FFC468", X"FFD972", X"FDDD6F", X"FFD262", X"FFCE65", X"F9CB6F", X"FDDA9D", X"705F55", X"0F0814", X"7A727C", X"F9F1F9"),
        (X"FEFFFF", X"7F828A", X"0E0E1B", X"615647", X"FADC8B", X"F8CF5D", X"FFD465", X"F9D363", X"F0D65F", X"FFDC77", X"F0AA6D", X"BE6141", X"D16756", X"C85D4D", X"BA5938", X"FDAF70", X"FFCB66", X"FAD05A", X"FCCF5C", X"F7D062", X"F4D76F", X"E1D287", X"4B4734", X"220F11", X"85493D", X"A95D37", X"C7863A", X"FFC75F", X"FFD75E", X"FBD459", X"FFDA6C", X"FFE085", X"FFE5A3", X"AE9C7E", X"221D2D", X"4D454E", X"E3CE9A", X"F5D87B", X"F7D968", X"EACD4C", X"EACF44", X"FFD758", X"FFB15A", X"B15620", X"AB5B3F", X"5E2614", X"311602", X"907B50", X"FFDF89", X"FCD364", X"F3D259", X"FAD75F", X"FFD763", X"FCCC61", X"C58C2B", X"A45A0D", X"B75522", X"BE4F2C", X"BC502E", X"BC4F30", X"BE4F30", X"BF593E", X"C06D59", X"804842", X"2E1C27", X"4C4538", X"F0D88A", X"F8D868", X"F4D461", X"F5D45F", X"FAD25D", X"FFCC5F", X"F7A246", X"B85601", X"C56A13", X"FFB75A", X"FFD56F", X"FFD467", X"F6D664", X"F7D863", X"FFD361", X"FFD067", X"FECA70", X"FFDA9E", X"705D54", X"130815", X"827781", X"FFFAFF"),
        (X"FEFFFF", X"7F8388", X"0E0E19", X"615645", X"FADD89", X"F8CF5D", X"FFD465", X"F9D363", X"F5DB64", X"F3D572", X"C29058", X"7C3A20", X"8C4038", X"86362D", X"863B20", X"DB9B63", X"FCCC6A", X"FAD05C", X"FCCF5C", X"F7D060", X"F2D56D", X"E2D389", X"494633", X"241115", X"854841", X"AA5D3F", X"C07D39", X"FFD171", X"FFD15C", X"FFD85E", X"FBD261", X"EECA67", X"E7CC78", X"A89563", X"2E2228", X"4D403D", X"E1C87E", X"F3D665", X"F5D661", X"F1D455", X"F0D44C", X"FCD058", X"FCAE60", X"BD6137", X"B66756", X"5A2318", X"2B1000", X"968156", X"FEDA84", X"FAD161", X"F3D058", X"F6D65D", X"F9D45F", X"FFD76A", X"E0AB49", X"CC8D37", X"E69853", X"E99659", X"E9955D", X"E89561", X"DD8C5C", X"9C5431", X"79442F", X"4F2D29", X"241923", X"464032", X"EAD284", X"F2D362", X"F4D461", X"F5D45F", X"FAD25D", X"FFCE5D", X"FCB24C", X"E59533", X"E29C34", X"FFC65B", X"FFCD5E", X"FCD462", X"F5D361", X"F0C95B", X"D99C38", X"DD973F", X"D89246", X"D9A371", X"5B433B", X"1B121E", X"7D727D", X"FFFDFF"),
        (X"FEFFFF", X"7F8386", X"0E0F13", X"61583D", X"FADD87", X"F8CF5D", X"FFD463", X"F9D363", X"F3D864", X"F7E081", X"AA935F", X"371C08", X"3C1F1B", X"3B1E1A", X"371901", X"C1A16C", X"F5D072", X"FCD15D", X"FDD05D", X"F8D261", X"EFD368", X"E4D48A", X"494535", X"25141A", X"854D47", X"BD7459", X"C07F43", X"FFC870", X"FFD76B", X"FFD15B", X"FDD05D", X"F3CB62", X"EFD678", X"AF995A", X"210800", X"4D321E", X"EBD079", X"F0D35F", X"F3D065", X"F3D063", X"F9DD62", X"FFD96E", X"F3AE6F", X"B9694B", X"AB6A62", X"623532", X"230F00", X"8E7E51", X"F6D981", X"F4D260", X"F4D55B", X"F5D65D", X"F7D35D", X"FDD165", X"FFCE6C", X"FFCD6F", X"FFD06A", X"FFD16D", X"FFD175", X"FFD17F", X"FED591", X"725528", X"261609", X"31292E", X"1B1827", X"443D30", X"E8D081", X"F0D060", X"F2D360", X"F4D25E", X"F9D05C", X"FAD05A", X"FCCF5A", X"FAD05A", X"F9D05C", X"F9D05C", X"FFD767", X"FAD066", X"FFDE79", X"E4A952", X"A9520F", X"B7501A", X"C05623", X"B2613F", X"533934", X"11101A", X"7D787E", X"FFFDFF"),
        (X"FEFFFF", X"7F8484", X"0E100F", X"615839", X"FADD87", X"F8CF5D", X"FFD463", X"F8D461", X"EFD75F", X"F1E381", X"9F9765", X"272214", X"29262C", X"282528", X"24210D", X"B4A574", X"F2D176", X"FCD05F", X"FDD05B", X"F8D25F", X"EDD166", X"E5D68B", X"484433", X"261622", X"78474E", X"905046", X"A4613A", X"F2B26F", X"F9BF63", X"FFD367", X"FED161", X"F9D466", X"F1D871", X"C2AD5D", X"63451D", X"6B4C1E", X"EED06F", X"F1D25D", X"F4CF65", X"F6CE67", X"F5CB61", X"F3C169", X"E2A16E", X"92543E", X"8D605D", X"523534", X"1B0E00", X"817748", X"F1D97F", X"F2D561", X"F4D85E", X"F6D85E", X"F8D45F", X"FDD165", X"FFCD6C", X"FFCC6A", X"FFD160", X"FFD25E", X"FFD167", X"FCD275", X"F3DB8F", X"655B2A", X"1B1B10", X"272D36", X"191B2A", X"453E31", X"E9D183", X"F1D161", X"F2D360", X"F4D25E", X"F9D05C", X"F7D25A", X"F2D45A", X"EFD55C", X"F1D45E", X"F2D360", X"FBD66A", X"FAD068", X"FFD878", X"F0B462", X"CC773B", X"DC7445", X"CB572C", X"BF6146", X"563734", X"111018", X"7C797E", X"FFFEFF"),
        (X"FEFFFF", X"7F8386", X"0E100F", X"61583B", X"FADD89", X"F8CF5F", X"FFD461", X"F8D55D", X"ECDA57", X"ECE77B", X"9A9967", X"22231A", X"242636", X"232633", X"212113", X"B1A776", X"F0D178", X"FCD05F", X"FDD05B", X"F8D25F", X"EDD164", X"E7D88B", X"494537", X"241A2E", X"32102B", X"400B1D", X"69241E", X"AF6442", X"B16A29", X"F8BC61", X"F5CC5F", X"FEE16D", X"E7D263", X"EAD574", X"E8CE7E", X"EBCD7C", X"F0CF64", X"F3D05A", X"F8CF5B", X"FECB5F", X"E7A449", X"A8611E", X"8C4E28", X"411403", X"402C2A", X"2B2522", X"211C0E", X"978E61", X"F0DA7F", X"F2D561", X"F3D95E", X"F4D85E", X"F8D45F", X"FDD165", X"FFCC6B", X"FFCA6A", X"FFCC61", X"FFCC5E", X"FFCA66", X"FACB72", X"F6DA8F", X"685A28", X"1E1A0B", X"2B2C34", X"191B2A", X"464032", X"E9D183", X"F2D362", X"F4D461", X"F5D45F", X"FAD25D", X"F8D25D", X"F2D35E", X"F1D460", X"F2D266", X"F6D068", X"F9D16D", X"F7CF6A", X"F9D36C", X"F3C769", X"FFC77B", X"FFBC7D", X"C9652E", X"BC6442", X"5B3530", X"180D16", X"7F797F", X"FFFFFF"),
        (X"FEFFFF", X"7F8386", X"0E100F", X"61583B", X"FADD89", X"F8CF5F", X"FFD461", X"F8D55B", X"EDDB59", X"EDE87C", X"9A996A", X"22231C", X"242638", X"232535", X"212115", X"B1A678", X"F0D178", X"FCD05F", X"FDD05B", X"F8D25D", X"EDD164", X"E7D88B", X"494537", X"211B30", X"321C3D", X"451C37", X"6A2932", X"A95C4B", X"AE632F", X"FFC574", X"F7D062", X"F7DD64", X"F6E06D", X"E7D062", X"E9CD63", X"EBCB5F", X"F8D461", X"F7CD57", X"FCCE57", X"FFC95F", X"E4934A", X"B56434", X"8E553B", X"3C1D13", X"252223", X"1B2524", X"181A0E", X"8E845C", X"F0DA82", X"F2D561", X"F2D85D", X"F2D65B", X"F8D45F", X"FDD165", X"FFCA6A", X"FFC66A", X"FFC267", X"FFC068", X"FFBF6B", X"FFC175", X"FED593", X"6D572C", X"22180E", X"2C2B34", X"1A1A2A", X"464032", X"E8D081", X"F2D362", X"F4D461", X"F5D45F", X"FAD25D", X"FCD15D", X"F9CF62", X"FACD68", X"FFCA6E", X"FFC872", X"FFC76F", X"FECB6C", X"F5CD64", X"F9D36C", X"F9CC72", X"FFCE7F", X"B96924", X"B87042", X"58372E", X"180B14", X"80787F", X"FFFDFF"),
        (X"FEFFFF", X"7F8386", X"0E100F", X"61583B", X"FADD89", X"F8CF5F", X"FFD461", X"F8D45F", X"F2DA65", X"F2E486", X"9C9368", X"1D1712", X"302D3C", X"2C2A36", X"2E281F", X"BCAC82", X"F1CF79", X"FACF5E", X"FCCF5A", X"F7D15C", X"EED363", X"E8D98C", X"4B4638", X"1F1E31", X"2E2739", X"391F2F", X"602B2F", X"A46050", X"AF6736", X"FDBF6D", X"FFDB66", X"F1D654", X"F4D860", X"F4D860", X"F7D85A", X"FBD658", X"FFD960", X"FDCB58", X"FFCA5B", X"FFCF74", X"E38B57", X"B15F46", X"88554B", X"2D1B1D", X"1C262E", X"16272D", X"181B16", X"8F855F", X"F3DD85", X"F2D561", X"EFD65A", X"EED358", X"F1CD58", X"FACE62", X"D49B3A", X"BC6E1E", X"D06726", X"D7622C", X"D2642E", X"C56936", X"B97D4D", X"5A3619", X"2D1F1F", X"33313F", X"1C1B2B", X"464032", X"E8D081", X"F4D463", X"F4D461", X"F5D45F", X"FAD25D", X"FFCE5F", X"F9B958", X"BE701F", X"C36928", X"C76A2C", X"B75E1A", X"EDA150", X"FFCF69", X"F8CA5F", X"FFD26F", X"FACC6E", X"F0BA63", X"F0C687", X"6B5C4A", X"110E13", X"827781", X"FFFBFF"),
        (X"FEFFFF", X"7E8486", X"0C110F", X"5F593B", X"F9DD89", X"F8CF5F", X"FFD461", X"F9D361", X"F7D769", X"F4DC82", X"9A8954", X"1D1100", X"221B0E", X"271F0F", X"1D1000", X"B5A168", X"F2CF74", X"FACF60", X"FCCF5A", X"F7D25A", X"EED363", X"E8D98C", X"4B4638", X"1F1E31", X"2F2C3B", X"2A1B27", X"542C35", X"9F6761", X"A76846", X"FCC07E", X"FFD46E", X"FFE16B", X"F7D662", X"F9D65E", X"FBD756", X"FFD755", X"FFD35B", X"FFCF60", X"FFC460", X"FFC77D", X"EB9B76", X"AD665C", X"845B5E", X"382A36", X"1E293A", X"1A2A37", X"1C1E1D", X"928867", X"F7E08B", X"F5D865", X"F2D85D", X"F0D459", X"FAD761", X"F7CB5F", X"C9902F", X"B26614", X"BC5418", X"C2501C", X"BE521C", X"B35722", X"A86A38", X"502B08", X"311E17", X"2A242C", X"1C1C29", X"464032", X"E6CF80", X"F5D565", X"F4D461", X"F5D45F", X"FAD25D", X"FFCD61", X"F9AC54", X"BF611D", X"C65A28", X"CB5A2E", X"C15822", X"F59D54", X"FFCE65", X"F8CC57", X"FFD96C", X"FED66D", X"F1CA68", X"F3D88F", X"655F48", X"0B0F12", X"7B7A81", X"FFFEFF"),
        (X"FEFFFF", X"7E8486", X"0C110F", X"5F593B", X"F9DD89", X"F8CF5F", X"FFD461", X"FDD25F", X"FACF60", X"FFDB76", X"D5BD68", X"96843B", X"9E904C", X"9D8F4B", X"A89449", X"E6CB75", X"F4D06A", X"FACF60", X"FCCF5A", X"F7D25A", X"EFD464", X"E9DB8E", X"4C473B", X"201F32", X"2A2738", X"281D2C", X"422639", X"6D444D", X"653027", X"C38966", X"C68E4D", X"EBB760", X"FCD26A", X"FCD462", X"FED45C", X"FFD35A", X"FFD158", X"FFD368", X"E7A251", X"DE9963", X"995B43", X"64332F", X"5F3C4A", X"34253C", X"1E233C", X"1B2337", X"1B181E", X"908365", X"F5DC87", X"F2D561", X"EED559", X"ECD056", X"F4D15B", X"FACE62", X"E9B04F", X"E8A64F", X"E29E4A", X"E49D4A", X"E59C4A", X"E19E4E", X"DAAC60", X"A9874C", X"A08C6C", X"6E645C", X"1D1C25", X"484133", X"E6CF80", X"F6D666", X"F5D563", X"F6D561", X"FBD35F", X"FFCE63", X"F7AC58", X"BF6023", X"C95730", X"CD5736", X"C25628", X"F39D56", X"FFD163", X"F2D053", X"FCDB62", X"FDDB6A", X"F7D168", X"FDE196", X"665F46", X"091010", X"708285", X"EFFFFF"),
        (X"FFFFFF", X"7E8488", X"0B0E14", X"615741", X"FEDA8F", X"FBCC65", X"FDD465", X"FBD261", X"FFD466", X"FFD369", X"F9D871", X"F8DD79", X"F7E07F", X"FCE584", X"F9DE7A", X"F8D971", X"F8D365", X"F9D05E", X"F9D15A", X"F7D15E", X"F4D166", X"F0D790", X"4F453B", X"221E34", X"242134", X"2B2338", X"312038", X"2C1023", X"380C10", X"9D6453", X"A35F34", X"DB9B56", X"FFD06E", X"FCD462", X"FFD35E", X"FFD25A", X"FFD256", X"FFD068", X"C87836", X"AA5F38", X"703E2F", X"37161B", X"3D273A", X"2C213E", X"242643", X"252840", X"201A23", X"99896E", X"FDE28E", X"FBDB66", X"F7DB60", X"F5D65D", X"FBD862", X"FFD86A", X"F9C561", X"FFCE6C", X"FFD26E", X"FFD36C", X"FFD16A", X"FFD16C", X"FBD172", X"F5D686", X"FAE6AD", X"9B8D70", X"201B1D", X"483F32", X"EBCC80", X"FBD464", X"F8D45F", X"F8D55D", X"F9D45D", X"FED067", X"F9B56D", X"BF6A39", X"C66148", X"CA624C", X"B75936", X"EA9F62", X"FDD36B", X"EDD255", X"F0D35B", X"F6D561", X"F5CE60", X"FEDF91", X"685F44", X"091010", X"708283", X"EDFFFF"),
        (X"FDFFFF", X"727781", X"0A091C", X"584441", X"E9B27E", X"EFB25B", X"F9CE68", X"FDDB6E", X"FBD265", X"F6CD60", X"F3CB60", X"F2CD63", X"F2CE66", X"F6D36B", X"F2CD63", X"F1CC5E", X"F2CF59", X"F3D058", X"F2D05C", X"F5CD62", X"EEBE5C", X"D8AE6F", X"57433C", X"262036", X"25213B", X"2A2640", X"2A213B", X"342133", X"4E292C", X"9A6253", X"B16541", X"F2A866", X"FFD56D", X"FDD961", X"FFD85D", X"FFD75B", X"FBD04F", X"FFD067", X"D7753D", X"BB5F48", X"764944", X"22131C", X"3B3348", X"24253E", X"20253F", X"2E2F43", X"1E1620", X"928066", X"F9DC86", X"F8D45F", X"F6D25C", X"F2CF59", X"FDD762", X"FAD15F", X"F8CD5E", X"F9CE5F", X"FAD161", X"FAD161", X"FFCF5D", X"FFCF5D", X"FFD669", X"EACA65", X"FCE892", X"978B54", X"211B16", X"4D3C32", X"F6CB83", X"FFD163", X"F9D053", X"F6D253", X"F3D357", X"F3CF6B", X"DEAD70", X"8F5234", X"8C443A", X"934B43", X"8C4B34", X"CF9A68", X"F9D67D", X"F8DD70", X"F5D565", X"F8D463", X"F5C958", X"FAD884", X"6B6248", X"0B0D0F", X"76787A", X"FDFFFF"),
        (X"FBFFFF", X"757B84", X"0E0A20", X"573D44", X"A86540", X"B66A26", X"F8C26B", X"FFD676", X"FFD16E", X"FFCC6A", X"FECA67", X"FFCB68", X"FFCC6A", X"FFD16E", X"FFCB68", X"FECA63", X"FECE5E", X"FFCE61", X"FFCD68", X"FFCA6E", X"AB6818", X"A97240", X"412926", X"251F35", X"272443", X"272445", X"272443", X"2F223B", X"3C1A25", X"97625B", X"B5674D", X"EB9D68", X"FFCA6E", X"FCCE60", X"FFCA5E", X"FFCA5C", X"FEC756", X"FFC96C", X"D27044", X"B45B50", X"70494B", X"221925", X"313247", X"242940", X"1D2239", X"212236", X"1B121E", X"9D8871", X"FFD989", X"FFD066", X"FFCE63", X"FBCB60", X"FFD469", X"FFCF65", X"FCCC61", X"FECD62", X"FFCF65", X"FFCF63", X"FFCE5F", X"FFCE5F", X"FFD367", X"FFD571", X"FFE68B", X"917F43", X"1D140E", X"523D34", X"F8C481", X"FFD26D", X"FFCF5D", X"FFD25B", X"FFD263", X"FCD179", X"D1A97B", X"421C0B", X"421B1A", X"3D1618", X"2F0800", X"A57D58", X"FBD28C", X"FFD57B", X"FED070", X"FFD16B", X"FCC75E", X"FFD788", X"665C44", X"0B0F12", X"7D7C7F", X"FFFDFF"),
        (X"F5FFFF", X"7A8085", X"140F21", X"56373F", X"AB6148", X"BB6230", X"FFAE6F", X"FFBE74", X"FFC171", X"FFBD6D", X"FFBA6A", X"FFBB6B", X"FFBD6D", X"FFC171", X"FFBB6B", X"FFBB66", X"FFBC63", X"FFBC65", X"FFB86B", X"FFB673", X"BE652C", X"B2714E", X"412A29", X"221E34", X"272447", X"27234B", X"27234B", X"2E2143", X"44273E", X"8A5961", X"985147", X"D78966", X"FFBA7A", X"FFBA6D", X"FFB66B", X"FFB569", X"FFB967", X"FFC17E", X"C47055", X"A25E5C", X"67494F", X"281F2B", X"2A2C40", X"262B42", X"1F243B", X"1F2034", X"221925", X"907565", X"FFCA89", X"FFBF68", X"FFBD65", X"FFB962", X"FFC26B", X"FFBE67", X"FFBA63", X"FFBB64", X"FFBE69", X"FFBE67", X"FFBC61", X"FFBC61", X"FFBF66", X"FFC271", X"FFCB84", X"A27E51", X"120201", X"523934", X"F0B07A", X"FFC777", X"FFC369", X"FFC367", X"FFC36B", X"FFC681", X"CBA486", X"35211C", X"322B2F", X"322A31", X"261512", X"A3806C", X"FFC698", X"FFC081", X"FFC276", X"FFC470", X"FFBC66", X"FFD08F", X"5C523E", X"0A1216", X"7D8688", X"FAFFFF"),
        (X"F2FFF8", X"7E8484", X"19131E", X"55343B", X"B56A5B", X"B95B39", X"C86438", X"C96432", X"CE6933", X"C9652C", X"C7632A", X"C8642B", X"C9652C", X"CE6A31", X"C8642B", X"C56428", X"C66625", X"CB6626", X"D3612A", X"D16032", X"BD5939", X"B36D5C", X"4D2E32", X"322A3F", X"292345", X"241F48", X"26214C", X"2F254B", X"37203C", X"4E2535", X"470A08", X"984E39", X"BC683E", X"C66632", X"D16030", X"D1612E", X"CD692F", X"CA7348", X"712A1D", X"4D1A20", X"624750", X"2C2430", X"2B2A3E", X"252A41", X"21273E", X"2D2C41", X"29202C", X"76534A", X"C47849", X"CD6A29", X"CA6827", X"C76424", X"D06D2D", X"CC6928", X"C86525", X"C86726", X"CA692A", X"CC6928", X"CF6822", X"CF6822", X"C76424", X"B86025", X"BA6D3E", X"814A2F", X"2E171A", X"4F302F", X"BA6E46", X"CF6E2F", X"CC6725", X"CE6723", X"CE6723", X"BF6A39", X"825544", X"221217", X"1A1C29", X"2B2F3E", X"2B1E25", X"7E544D", X"C36C53", X"C86036", X"C9652E", X"C76929", X"BC6020", X"B97648", X"5C463E", X"0E121A", X"82888F", X"FAFFFF"),
        (X"F6FFF5", X"757A74", X"090207", X"44262C", X"B06D66", X"BB604F", X"C0573D", X"C24C30", X"D65A3B", X"D55434", X"D35132", X"D45333", X"D55434", X"DA5839", X"D45333", X"CF5332", X"CA582F", X"CB5930", X"D35532", X"CF553C", X"C36056", X"A85E60", X"421922", X"2B1628", X"271B36", X"211B3D", X"232247", X"302D4E", X"3A2A46", X"3C1E2F", X"451719", X"864438", X"B95D45", X"C7573B", X"CD5539", X"CD5537", X"CA5D37", X"BC6348", X"632A2B", X"371523", X"4E3844", X"312635", X"2D2C3F", X"25283E", X"202439", X"252437", X"2D2131", X"714645", X"C05E43", X"D05029", X"D3532C", X"D3532C", X"D3532C", X"D1512B", X"D3532C", X"D35530", X"D15531", X"D1532E", X"D65228", X"D65228", X"D5552E", X"C65031", X"C85E49", X"8C3D36", X"3A1620", X"532C30", X"B45F45", X"C75B32", X"C9592F", X"CA592D", X"CA592B", X"BC5D3D", X"925855", X"381A2B", X"262036", X"29253D", X"351C2D", X"85464E", X"CF5D53", X"DE553F", X"D35230", X"CE552E", X"CB5630", X"B65D44", X"60393B", X"201424", X"787483", X"FFFDFF"),
        (X"FBFFF2", X"D1D6C9", X"B5AEAC", X"9B8283", X"693535", X"80312C", X"BF5A4E", X"CA5646", X"D45545", X"D34F40", X"D04C3E", X"D14D3F", X"D34F40", X"D75345", X"D14D3F", X"CD4E3C", X"C8533B", X"C7553C", X"CC533A", X"C45546", X"80292D", X"74303E", X"7A4353", X"714A5B", X"362536", X"232033", X"22253D", X"30334B", X"342E42", X"34222D", X"3D1B19", X"81463A", X"BC5F4F", X"CA5947", X"CC5945", X"CC5943", X"C15739", X"B55F4C", X"5B2D33", X"32182A", X"493744", X"362B3A", X"2C2B3E", X"25283E", X"1F2338", X"252437", X"2D2131", X"714549", X"C55E51", X"D4513B", X"D6533D", X"D6533D", X"D6533D", X"D5523C", X"D6533D", X"D85640", X"D65541", X"D6533D", X"DB5237", X"DB5237", X"D8563E", X"CB5041", X"CD5F59", X"913E43", X"431826", X"592C34", X"B45B4E", X"C4533C", X"C2523A", X"C25238", X"C15434", X"B45841", X"8E5254", X"39182A", X"2A2139", X"312842", X"321629", X"8C4D55", X"D35E56", X"D04633", X"D6543B", X"D1563D", X"CE5741", X"B95E54", X"684047", X"180C1E", X"7C7489", X"FFF9FF"),
        (X"FFFFF4", X"FFFFFB", X"FFFEF6", X"C5B6B4", X"270507", X"4C1515", X"A95852", X"CA675D", X"CE6257", X"CC5C52", X"CA5A50", X"CB5B51", X"CC5C52", X"D16157", X"CB5B51", X"C85B4E", X"C85D4F", X"C85F4E", X"C6614C", X"BB6458", X"41020E", X"50162C", X"A1596F", X"AD7181", X"4A3238", X"2C2C2E", X"242C32", X"2C333C", X"2E3137", X"2E2725", X"372011", X"7B4A36", X"B96350", X"C45E4A", X"C06146", X"BF6244", X"C76A4A", X"B86B58", X"5A3136", X"2E1728", X"473541", X"3C3040", X"252437", X"272B3E", X"1F2336", X"252437", X"2D2131", X"6E464B", X"B9645A", X"C55846", X"C85C4A", X"C75B49", X"C75B49", X"C65948", X"C75B49", X"CA5D4D", X"C75C4C", X"C75B49", X"CC5943", X"CC5943", X"CB5D49", X"BE574C", X"BE6664", X"88434A", X"390D1E", X"592432", X"BB5E59", X"CB5D50", X"C55E53", X"C06151", X"BD6449", X"B06951", X"8F625C", X"392129", X"231F2E", X"231E30", X"2F1B24", X"7E4D47", X"C56C53", X"D36747", X"CB5F46", X"C8604A", X"C66050", X"B36660", X"51343C", X"0C091A", X"6C6A82", X"FEFFFF"),
        (X"FEFFF2", X"FDFDEF", X"FCFBF2", X"D9D0CF", X"7E6B6D", X"825F62", X"864F4D", X"8B4745", X"914946", X"8E4441", X"8C413F", X"8D4240", X"8E4441", X"934846", X"8D4240", X"8C4141", X"8F4144", X"8E4343", X"8D453D", X"884643", X"6A2E40", X"6F304A", X"843B54", X"844452", X"5B3A37", X"3E3027", X"2D2B29", X"2F3133", X"302F32", X"2C2827", X"2F221B", X"6E4D44", X"884A3F", X"8F4739", X"8B4939", X"894A39", X"854431", X"8B5248", X"4F2934", X"351E2E", X"443241", X"3F3443", X"252233", X"2A2D41", X"1F2336", X"282536", X"2D2131", X"664953", X"854C4D", X"89433F", X"8B4541", X"8B4541", X"8B4541", X"8A4440", X"8B4541", X"8D4744", X"8E4641", X"8E443D", X"92433B", X"92433B", X"924640", X"883F3F", X"8F4B55", X"612633", X"5B2D3D", X"65313E", X"9E545B", X"944348", X"8E4449", X"894747", X"864A3F", X"7E4E41", X"664643", X"291419", X"3A2833", X"4F3B44", X"55373A", X"673C36", X"834634", X"944E38", X"8C4634", X"8C4538", X"8C443C", X"7D4946", X"6C5B61", X"686A77", X"9C9EB0", X"FEFFFF"),
        (X"FDFBF9", X"FEFCFB", X"FEFCFB", X"FFFBFD", X"FFFFFF", X"FFF4F6", X"3E2B2D", X"2B1317", X"311823", X"321828", X"2D1423", X"341B2A", X"3C2332", X"391F2F", X"341B2A", X"32182A", X"341731", X"3A1B31", X"3C1F27", X"461922", X"AE6479", X"B06179", X"450A20", X"410F1B", X"925F59", X"9A6E64", X"513636", X"3A292F", X"372831", X"493D4C", X"524C62", X"2A2033", X"3A2228", X"3D2124", X"38232A", X"37232E", X"341A25", X"371A28", X"674757", X"3D2131", X"342030", X"4E4050", X"292637", X"242638", X"27283A", X"282536", X"372939", X"4A394A", X"2E2033", X"2E2035", X"2E2035", X"2E2035", X"2E2035", X"2D1E33", X"2E2035", X"322233", X"34212A", X"361E28", X"381C2E", X"3A1B31", X"331828", X"371628", X"360922", X"522136", X"986771", X"8E626A", X"39182A", X"2D1329", X"31162D", X"2C1226", X"2F1A26", X"301C25", X"26151D", X"32181F", X"815259", X"A87075", X"A87075", X"65363D", X"341721", X"301C25", X"311A1B", X"2C1313", X"331A1C", X"1D0A0E", X"BFB9BF", X"F9FAFF", X"FDFEFF", X"FBFCFF"),
        (X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FFFFFF", X"EEEBEE", X"474749", X"3D3B43", X"424252", X"302F44", X"2A2C40", X"313247", X"222337", X"26273B", X"2A2C40", X"2D2B43", X"2B2645", X"292240", X"282335", X"351E2C", X"8E4F64", X"853B52", X"6C3246", X"5D2730", X"995F5A", X"A3695F", X"582B28", X"4B282D", X"3B2432", X"4A3B52", X"524A6B", X"25213D", X"2C2734", X"2C2832", X"27283C", X"272740", X"261F3A", X"2C1C36", X"5C4053", X"432536", X"3B2334", X"483A4A", X"292637", X"262739", X"232537", X"232031", X"3E2F42", X"493F53", X"20253F", X"1B2645", X"1B2645", X"1B2645", X"1B2645", X"1A2544", X"1B2645", X"1F2943", X"23263A", X"232539", X"232343", X"252145", X"221D3C", X"3A2843", X"452035", X"663646", X"85565F", X"775561", X"32283C", X"272541", X"2A2341", X"382C49", X"2C2334", X"291A23", X"391A20", X"4B1F22", X"783E44", X"8F525B", X"85515E", X"553446", X"282237", X"262C3E", X"34353E", X"3B3B3F", X"46454A", X"38373C", X"BEBDC4", X"FDFCFF", X"FAFAFC", X"FFFFFF"),
        (X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"F8F5FB", X"FDFAFF", X"FCFBFF", X"F3F2F9", X"FAFAFF", X"8A8A98", X"1D202D", X"212330", X"1A1C2B", X"1D1F2F", X"222433", X"262636", X"292438", X"262339", X"24253C", X"29233A", X"280E25", X"431227", X"A85F71", X"B86B75", X"632825", X"58231A", X"9C6258", X"9A6867", X"3D2133", X"4A3B55", X"584960", X"2C2031", X"2F2630", X"2C2832", X"28273C", X"282640", X"28213D", X"2D1E37", X"523648", X"4A2C3D", X"2B1425", X"3F3141", X"2A2836", X"3D3F4E", X"3B3D4C", X"252233", X"3B2C41", X"34273E", X"22253B", X"1D273F", X"1D2641", X"1D2641", X"1D2641", X"1C253F", X"1D2641", X"212843", X"242540", X"23233F", X"202541", X"222343", X"2D2449", X"3C2340", X"996870", X"946062", X"391223", X"361E32", X"2E2330", X"352B3C", X"35223F", X"361D38", X"341A21", X"7A524B", X"B36E63", X"A45C57", X"66303B", X"3A172E", X"261632", X"26243C", X"1F2631", X"11191F", X"727379", X"F5F4F9", X"F0EFF4", X"F7F6FB", X"F8F7FC", X"FFFFFF", X"F7F6F9", X"FFFFFF"),
        (X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"F5F2F7", X"FFFFFF", X"FEFDFF", X"FDFBFF", X"FDFFFF", X"A3A3AC", X"3D4048", X"4F535B", X"343641", X"31343E", X"2D2F3A", X"292A35", X"2C2535", X"2B2338", X"29223E", X"292240", X"2E283E", X"3F2535", X"955863", X"A15A5E", X"632D26", X"542218", X"975B52", X"A46C6A", X"461D2B", X"56374A", X"5F4856", X"2F2029", X"2F272E", X"2C2832", X"28273C", X"282640", X"2A243F", X"2E1F39", X"492D40", X"503243", X"382132", X"473949", X"27222F", X"2E303D", X"363845", X"201B2C", X"423348", X"392A3F", X"252439", X"20263B", X"20263B", X"20253D", X"20253D", X"1F243B", X"20253D", X"242641", X"262342", X"252241", X"22253D", X"26223B", X"3F2844", X"4C273A", X"916162", X"7D504F", X"3B2133", X"2C1F33", X"28222B", X"271B23", X"48273B", X"5C3041", X"461A1B", X"804A45", X"A25853", X"A25C5D", X"592E3F", X"2F1B34", X"292A40", X"414A59", X"454F4E", X"2E332F", X"8C8B8E", X"FEFDFF", X"FFFFFF", X"FAFAFE", X"FFFEFF", X"FCFBFF", X"FFFFFF", X"FFFFFF"),
        (X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FDFCFF", X"FDFCFF", X"FBFDFF", X"FBFCFF", X"FBFCFF", X"FBFCFF", X"E3E4EA", X"26272E", X"191C22", X"25242D", X"1B1220", X"35213A", X"3A183D", X"2C0F34", X"2A243B", X"2A272F", X"372321", X"412015", X"896151", X"946459", X"80494C", X"5C1F26", X"AC6C6D", X"875051", X"422427", X"66575C", X"544C51", X"27232D", X"2B2A3E", X"1F1D37", X"1C1631", X"2D1E37", X"3B1F32", X"593B4C", X"351E2E", X"473748", X"342F3C", X"20212C", X"1D1D2A", X"211C2C", X"4B3A4D", X"3A293F", X"292436", X"262538", X"262538", X"252437", X"212133", X"1F1E31", X"201F32", X"25233B", X"251F44", X"292345", X"2C253E", X"402C39", X"956268", X"915B5B", X"452021", X"321D22", X"28242C", X"1B1E28", X"232631", X"2A1B23", X"885154", X"AE676A", X"A16068", X"662D3C", X"48162E", X"401932", X"33192D", X"20131F", X"494448", X"FEFDF7", X"FCFCEE", X"F8F5E8", X"FFFBFB", X"FEFBFF", X"FDFCFF", X"FDFCFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF"),
        (X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FEFBFF", X"FDFCFF", X"FDFCFF", X"FBFDFF", X"FBFDFF", X"FBFDFF", X"FBFDFF", X"F3F5F7", X"636566", X"4D5252", X"2D2E35", X"362F41", X"34203B", X"462044", X"462645", X"383443", X"34383B", X"383731", X"403529", X"806352", X"906458", X"7D4347", X"551218", X"B26360", X"B36D67", X"3F1914", X"73625E", X"60565A", X"27232D", X"2E2D42", X"33314B", X"352E49", X"43344E", X"4D3143", X"6A495B", X"3D2435", X"3D2C3D", X"2A2631", X"82838C", X"747480", X"201B2A", X"4D3C50", X"48384B", X"3E3445", X"3B3547", X"3B3547", X"3B3645", X"383443", X"373242", X"383443", X"3F374C", X"3F3352", X"3A2847", X"3C2437", X"4B282F", X"9F6663", X"915C55", X"4B2F32", X"34282E", X"353034", X"3D353A", X"3E2A31", X"421F22", X"8C554C", X"9C5E58", X"8D535D", X"5B2C43", X"462849", X"3E2D4C", X"403747", X"575055", X"767069", X"FFFBED", X"FFFBEB", X"FFFFFF", X"FFFBFB", X"FEFBFF", X"FDFCFF", X"FDFCFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF"),
        (X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FEFEFE", X"FEFEFE", X"FCFFFE", X"FCFFFE", X"FCFFFC", X"FCFFFC", X"FFFFFE", X"F6F9F6", X"F9FFFB", X"EAEEF4", X"8E8CA3", X"241A39", X"342037", X"3E2C39", X"322D2F", X"302E2D", X"322D2F", X"372B2B", X"3C271C", X"451B10", X"722F2A", X"A95758", X"9C4A4B", X"97514D", X"75483A", X"856C60", X"382C2C", X"908C96", X"9E9BB0", X"15112B", X"29223E", X"34253E", X"391D30", X"513143", X"4B3243", X"342332", X"1E1A24", X"A8A9B2", X"B9BAC2", X"25202D", X"4F3F50", X"342133", X"2E2232", X"2C2334", X"2C2334", X"2E2433", X"2E2433", X"2E2433", X"2F2634", X"372939", X"472C43", X"4A243A", X"7C4B57", X"8E5B61", X"3F1918", X"412422", X"3C262B", X"432D32", X"422429", X"845457", X"A15656", X"AC645F", X"492417", X"3F2C25", X"3D252D", X"331E31", X"201129", X"BCB6CA", X"FFFFFF", X"FDFFFE", X"FCFDF3", X"FFFCF3", X"FFFFFB", X"FFFBFA", X"FFFBFE", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF"),
        (X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FFFDFF", X"FEFEFE", X"FEFEFE", X"FCFFFC", X"FCFFFC", X"FCFFFC", X"FCFFFC", X"FFFFFF", X"FFFFFF", X"F6FBF7", X"FEFFFF", X"B4B5C9", X"5B576F", X"564F5B", X"2B2426", X"403C39", X"403C39", X"403B3F", X"43393F", X"4E3A3A", X"582F2D", X"833F3C", X"B46262", X"9C4C4C", X"490100", X"C08874", X"AE8875", X"342423", X"A19DA8", X"B3B1C1", X"171429", X"403B51", X"483B4F", X"473041", X"5C4350", X"4D3645", X"3F2F3E", X"45424A", X"C8C9CF", X"ACADB4", X"1C1823", X"554554", X"443241", X"473443", X"453545", X"453545", X"463645", X"4A3A48", X"4A3A48", X"4B3B49", X"563D4C", X"43192A", X"511C29", X"8F5960", X"815559", X"50393A", X"422F34", X"44262C", X"42181F", X"57212A", X"9C575E", X"C36869", X"B66B67", X"574036", X"32332C", X"383238", X"635C6A", X"5E5765", X"DAD8E2", X"F1F6F7", X"F6FDF8", X"F4F8F0", X"FEFAF2", X"FFF8F7", X"FFF9FA", X"FFFCFE", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF", X"FEFDFF"),
        (X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FCFFFE", X"FCFFFE", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FCFDFF", X"FFFFFF", X"F5F2F5", X"CDCBCC", X"3B3937", X"252221", X"3E3C3D", X"433941", X"4A3140", X"522939", X"58202C", X"5B1B1E", X"611B18", X"A05749", X"A45A43", X"A56D59", X"463230", X"939098", X"F8F6FF", X"B9B7C3", X"373340", X"342E39", X"3A2F39", X"3B2E37", X"55424F", X"382A36", X"CBC7CF", X"FFFFFF", X"AAABB1", X"1F1B23", X"423540", X"3E2937", X"442B3A", X"462A3C", X"462A3C", X"462A3C", X"3D2133", X"44283A", X"482C3F", X"4D2537", X"7F414F", X"90535C", X"432025", X"433135", X"473B3F", X"493137", X"804A51", X"9B555F", X"934A5C", X"651E30", X"61222B", X"42171A", X"261615", X"898783", X"E2E0E1", X"FFFDFF", X"FFFCFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFFFC", X"FEFDF9", X"FFFDFB", X"FFFDFD", X"FFFDFE", X"FEFDFF", X"FFFDFF", X"FFFDFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FCFFFE", X"FCFFFE", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FCFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"808080", X"717171", X"2F2F2F", X"362E35", X"5A4055", X"613B53", X"623949", X"663740", X"7E4745", X"B47B6E", X"A56652", X"410F00", X"BBA9A9", X"F6F3FB", X"FFFFFF", X"F3F2F9", X"1C1921", X"39363E", X"4A474C", X"504850", X"675763", X"261924", X"CAC6CE", X"FAFBFF", X"9FA1A5", X"1B181E", X"655861", X"4E3A45", X"5B3F4F", X"5D3E4F", X"5D3E4F", X"5D3E4F", X"5F4054", X"5B3D50", X"3A1B2E", X"2D0616", X"985D66", X"9C696F", X"564548", X"373639", X"111113", X"29191C", X"925F65", X"B16D76", X"AE6C7B", X"6D3445", X"38121C", X"7E696E", X"6C6263", X"C1BFBD", X"FFFFFF", X"F8F6F5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFFFFD", X"FFFFFD", X"FFFFFD", X"FFFEFF", X"FEFDFF", X"FEFDFF", X"FFFDFF", X"FFFDFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFBFC", X"FAFAFA", X"FEFEFE", X"F9F9F9", X"FFFFFF", X"D5D5D7", X"7A747B", X"402E3A", X"462C3E", X"492E3C", X"4C313C", X"45292E", X"422627", X"4A2F2B", X"B4A09D", X"F5EBEF", X"FFFFFF", X"FFFEFF", X"F3F2F9", X"C3BFC7", X"49454D", X"2F2C31", X"3C333B", X"43333D", X"C3B7BF", X"F1EEF6", X"FFFFFF", X"E6E8EC", X"A3A1A4", X"42353E", X"422E3A", X"4A313E", X"4C303E", X"4C3040", X"4C3040", X"4B2F3F", X"3A1F2F", X"836679", X"AD8F9E", X"3C1E24", X"3B2425", X"343132", X"6C7373", X"B8BFBF", X"A5A2A3", X"4D3636", X"442126", X"442128", X"705459", X"C5B7B9", X"FBF7F6", X"FDFDFB", X"FBFEFB", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFFBFB", X"FFFDFC", X"FFFDFC", X"FFFDFC", X"FFFFFD", X"FFFEFF", X"FFFEFF", X"FFFEFF", X"FFFEFF", X"FFFEFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FDFFFF", X"FFFFFF", X"FFFFFF", X"F7F7F7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFBFC", X"FDFDFD", X"FDFCFF", X"CAC5CB", X"7D6D79", X"846F7D", X"877581", X"8B7986", X"8D7E88", X"8A7E84", X"8D8487", X"FFFEFF", X"FFFDFF", X"FAF6FC", X"F8F7FE", X"FFFFFF", X"FFFFFF", X"928E96", X"7A767C", X"7D757C", X"8F808A", X"FFFEFF", X"FEFBFF", X"FFFFFF", X"F6F8FC", X"F4F1F4", X"867982", X"8E7A85", X"8A737F", X"8B737F", X"8B7281", X"8B7281", X"8D7383", X"89707F", X"CBB2C4", X"FCE5F2", X"927F83", X"857C7B", X"686D6B", X"BECAC8", X"F7FFFF", X"FCFFFF", X"8F8586", X"857274", X"836E70", X"AE9E9F", X"FFFFFF", X"FBFEFB", X"FCFFFD", X"FAFDF9", X"FCF8F7", X"FFF6F7", X"FFF8F8", X"FFFBFB", X"FFFBFB", X"FFFDFC", X"FFFDFC", X"FFFDFC", X"FFFFFD", X"FFFEFF", X"FFFEFF", X"FFFEFF", X"FFFEFF", X"FFFEFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF")
    );

    
    constant win: winArray := (
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"FFF9BD", X"FFF9BD", X"FFC20E", X"FFC20E", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"FFC20E", X"FFC20E", X"FFF9BD", X"FFC20E", X"FFC20E", X"FFC20E", X"D4BB00", X"FFC20E", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"FFFFFF", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"D4BB00", X"FFFFFF", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"FFC20E", X"D4BB00", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"FFC20E", X"FFC20E", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFC20E", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"000000", X"000000", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"D4BB00", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"D4BB00", X"D4BB00", X"D4BB00", X"D4BB00", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF")
    );

    constant AFLOGO: LOGOArray := (
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF4F7", X"FDE5EB", X"FEF6F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FDFDFD", X"FDFDFD", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDFE7", X"F47E9D", X"F1577F", X"F47F9D", X"FCDCE4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FBFBFB", X"F8F8F8", X"F7F7F7", X"F6F6F6", X"F6F6F6", X"F7F7F7", X"FAFAFA", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDE6EC", X"F37092", X"EF406D", X"EF406E", X"EF3F6D", X"F37394", X"FDEBF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFD", X"F697B0", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF4471", X"F7A5BA", X"FFFEFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDFE7", X"F15A81", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F26086", X"FDE2E9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F6F6F6", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8A9BD", X"EF4370", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4370", X"F8AABE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FCFCFC", X"FEFEFE", X"FDFDFD", X"FBFBFB", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF6F8", X"F47A99", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F47A99", X"FEF6F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCE1E8", X"F1587F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F1577F", X"FDE0E7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC3D2", X"F04975", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"F04974", X"FAC0CF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F7A3B9", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F8A4BA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"F58AA6", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F691AC", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF4F6", X"F37394", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F482A0", X"FEF9FA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEEFF3", X"F26489", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F37797", X"FEF5F7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDECF1", X"F15C83", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F36F91", X"FEF2F5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF1F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FDFDFD", X"FEFEFE", X"FEFEFE", X"FCFCFC", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F6F6F6", X"F6F6F6", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF6F9", X"FAC0CF", X"FCDCE4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"FBCBD8", X"FBCBD7", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFE", X"F8A8BD", X"EF4773", X"F2698D", X"FDE3EA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBCAD6", X"F0537C", X"F0527B", X"FAC7D4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FBFBFB", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDCE4", X"F15B82", X"EF406D", X"EF426F", X"F699B1", X"FFFCFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8F9", X"F5829F", X"EF3F6D", X"EF406D", X"F37697", X"FEF1F5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FBFBFB", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F8F8F8", X"F7F7F7", X"F6F6F6", X"F6F6F6", X"F8F8F8", X"FAFAFA", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8B1C3", X"EF4370", X"EF426F", X"EF406E", X"F26187", X"FDEAEF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDFE7", X"F1567E", X"EF416E", X"EF416E", X"F04D77", X"FBCCD8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFD", X"F68FAA", X"EF3F6D", X"EF426F", X"EF416E", X"F04B76", X"FAC9D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9B9CA", X"EF4672", X"EF426F", X"EF426F", X"EF416F", X"F7A5BB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF4F7", X"F37596", X"EF406D", X"EF426F", X"EF426F", X"EF4470", X"F8B0C3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEDF1", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F2698D", X"FEF3F6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F79AB2", X"EF3F6D", X"EF426F", X"EF426F", X"EF3F6D", X"F58BA7", X"FFFCFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEEFF3", X"F26489", X"EF406E", X"EF426F", X"EF426F", X"EF416E", X"F7A7BC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFD", X"FDE6EC", X"FAC4D2", X"FABECE", X"FABECE", X"FABECE", X"FABFCF", X"F8B1C4", X"F05079", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F26186", X"F9B6C8", X"FABFCE", X"FABECE", X"FABECE", X"F9BECD", X"FBCDD9", X"FEF2F5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"F589A5", X"EF3F6D", X"EF426F", X"EF426F", X"EF3F6D", X"F482A0", X"FEF9FA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBF0", X"F1587F", X"EF416E", X"EF426F", X"EF426F", X"EF3F6C", X"F7A1B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEEFF3", X"FAC6D4", X"F690AA", X"F15E85", X"F04975", X"EF4773", X"EF4773", X"EF4773", X"EF4773", X"EF4672", X"EF436F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4572", X"EF4773", X"EF4773", X"EF4773", X"EF4773", X"EF4773", X"F04D78", X"F36E90", X"F7A5BB", X"FCD8E2", X"FEF8F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF7F9", X"F47C9B", X"EF3F6D", X"EF426F", X"EF426F", X"EF3F6D", X"F47C9B", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF6F8", X"FBD4DE", X"F7A1B7", X"F26A8D", X"F04B75", X"EF406D", X"EF406E", X"EF416E", X"EF416F", X"EF416F", X"EF416F", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"EF416F", X"EF416F", X"EF416F", X"EF426F", X"EF416E", X"EF406D", X"EF426F", X"F0547C", X"F47D9C", X"F8B4C6", X"FDE4EA", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF6F8", X"F37B9A", X"EF406D", X"EF426F", X"EF426F", X"EF406D", X"F37B9A", X"FEF6F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF3E6C", X"F7A1B8", X"FFFFFF", X"FFFBFC", X"FCE1E8", X"F8B0C2", X"F47999", X"F0517B", X"EF416E", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF3F6D", X"EF4571", X"F15C83", X"F58BA7", X"FAC2D1", X"FDECF0", X"FFFFFF", X"FEF9FA", X"F47C9B", X"EF3F6D", X"EF426F", X"EF426F", X"EF406D", X"F37B9A", X"FEF6F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF3F6D", X"F691AB", X"FAC5D3", X"F589A5", X"F15A81", X"EF4471", X"EF3F6D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"EF406D", X"F04974", X"F2678B", X"F699B1", X"FAC6D4", X"F37696", X"EF406D", X"EF426F", X"EF426F", X"EF406D", X"F37B9A", X"FEF6F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBF0", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"F04D77", X"F04A75", X"EF406D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF406E", X"F04E78", X"F04C76", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F37C9B", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDE6EC", X"F1557E", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F37898", X"FEF4F6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFD", X"FDE6EC", X"F9B8C9", X"F47B9A", X"EF4672", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"F04E78", X"F58BA7", X"FAC4D2", X"FEF0F3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF0F3", X"FAC5D3", X"F68FA9", X"F15D83", X"EF4571", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"F04975", X"F2698D", X"F7A0B7", X"FCD5DF", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"FBFBFB", X"FAFAFA", X"FBFBFB", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"F9F9F9", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF6F8", X"FBD4DE", X"F7A0B6", X"F2698C", X"F04A75", X"EF3F6D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF406E", X"F0517A", X"F37797", X"F8B1C4", X"FDE2E9", X"FFFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"FDE1E8", X"F8AFC2", X"F37697", X"F0517A", X"EF406E", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF4370", X"F15A81", X"F58AA5", X"FAC1D0", X"FDEDF1", X"FFFEFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFE", X"FDEBF0", X"FABFCE", X"F587A3", X"F15981", X"EF4370", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"EF3F6D", X"F04873", X"F2668A", X"F79BB3", X"FBD1DC", X"FEF5F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F7F7F7", X"FAFAFA", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF4F7", X"FBCEDA", X"F698B0", X"F26489", X"EF4773", X"EF3F6D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"EF406D", X"EF406E", X"F04F79", X"F37395", X"F8ACC0", X"FCDEE6", X"FFFAFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"F9F9F9", X"FAFAFA", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FBFBFB", X"FBFBFB", X"FCFCFC", X"FDFDFD", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9FB", X"FCDBE4", X"F8A9BE", X"F37193", X"F04E78", X"EF406E", X"EF406D", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF426F", X"F15880", X"F584A1", X"F9BCCC", X"FDEAEF", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFE", X"FDE8ED", X"F9B9C9", X"F4819F", X"F1567E", X"EF426F", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"EF3F6D", X"EF4773", X"F26288", X"F696AF", X"FBCCD8", X"FEF2F5", X"FFFFFF", X"FDFEFE", X"F6F7F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF0F4", X"FAC9D6", X"F692AC", X"F26186", X"EF4672", X"EF3F6D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"EF406E", X"F04D77", X"F37092", X"F6A5BA", X"F4D3DB", X"F4EFF0", X"F5F7F6", X"F5F7F6", X"F9FAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"FCD7E1", X"F7A4BA", X"F36D90", X"F04C76", X"EF406E", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EA406C", X"E75179", X"EB7997", X"EFAFC0", X"F6DEE4", X"FEFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFD", X"FDE4EA", X"F9B4C6", X"F47D9C", X"F0547C", X"EF426F", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426E", X"E73F6B", X"E63E6A", X"E63D69", X"E7436E", X"EF5C82", X"F68EA9", X"FAC6D3", X"FEEEF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEEEF2", X"FAC6D4", X"F58EA9", X"F15D84", X"EF4571", X"EF3F6D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EC416D", X"E63F6B", X"E63F6B", X"E63F6B", X"E83F6C", X"EE406D", X"EF406D", X"F04A75", X"F36A8E", X"F79EB5", X"FBD3DD", X"FEF5F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9FB", X"FBD4DF", X"F79FB6", X"F36B8E", X"F04A75", X"EF406D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EA406D", X"E63F6B", X"E63F6B", X"E63F6B", X"EA406D", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF416E", X"F0517B", X"F37798", X"F8AFC2", X"FCE0E7", X"FFFDFD", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDFE6", X"F588A4", X"F0537C", X"EF416E", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"E9406D", X"E63F6B", X"E63F6B", X"E63F6B", X"E9406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF4470", X"F15B82", X"F7A1B8", X"FBECF0", X"F6F7F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEDF1", X"F37193", X"EF3F6D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EA406D", X"E63F6B", X"E63F6B", X"E63F6B", X"E8406C", X"EE426E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"ED436F", X"EE8BA5", X"F4EFF1", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FACAD6", X"F04B75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EB416D", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"EA406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"ED416E", X"E83E6A", X"E8567D", X"F3E3E7", X"F5F6F6", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCD8E1", X"F1547D", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426E", X"E73F6C", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"EA416D", X"EE426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"EB416D", X"E73F6B", X"E63C69", X"EA6D8E", X"F4E9EC", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"F8A8BD", X"F1557E", X"EF4370", X"EF406D", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF3F6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EA3D6A", X"E63B68", X"E63B68", X"E63B68", X"E63B68", X"E63C68", X"E83C69", X"EA3D6A", X"EB3D6B", X"E93D6A", X"E73C69", X"E63E6B", X"E6436E", X"E96688", X"F1C7D2", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFC", X"FCD9E2", X"F8ACC0", X"F694AD", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F4809E", X"F04A75", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F0507A", X"F482A0", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F487A4", X"EE85A0", X"EB829E", X"EC829E", X"EC829E", X"EC829E", X"EB829E", X"EB829E", X"EB829E", X"EB829E", X"EC85A0", X"ED97AD", X"EFB4C4", X"F4E1E6", X"F9FAF9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDECF0", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF2F5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFFFF", X"F8FAF9", X"F5F7F6", X"F5F6F6", X"F5F7F6", X"F5F7F6", X"F5F7F6", X"F5F7F6", X"F5F7F6", X"F5F6F6", X"F5F7F6", X"F7F9F8", X"FBFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"FAFAFA", X"F9F9F9", X"FBFBFB", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F9F9F9", X"F6F6F6", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FDFDFD", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FBFBFB", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEAEF", X"F1577F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2698D", X"FEF0F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F7F7F7", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBF0", X"F1567F", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F26A8D", X"FEF3F6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"FCD7E0", X"F79EB5", X"F04A75", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F15B82", X"F9B8C9", X"FDEAEF", X"FFFEFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFD", X"FDE1E8", X"F9B2C5", X"F47999", X"F0527B", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4672", X"F26388", X"F694AE", X"F9CBD7", X"F8EDF0", X"FDFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBEF", X"F9C0CF", X"F586A3", X"F15A81", X"EF436F", X"EF3F6D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"EC3F6C", X"E84973", X"E9688A", X"F09FB5", X"FBD7E0", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF2F5", X"FBCFDA", X"F697AF", X"F26489", X"EF4773", X"EF406D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EC416E", X"E73F6B", X"E63E6A", X"E63D69", X"E63E6A", X"EB5179", X"F37999", X"F8B1C3", X"FCE1E8", X"FFFBFC", X"FEFFFF", X"F7F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FBFBFB", X"FAFAFA", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF9FA", X"FCDBE3", X"F7A7BC", X"F37293", X"F04D77", X"EF406E", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EC416E", X"E73F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63E6A", X"EA3E6B", X"EF4370", X"F15A81", X"F585A2", X"F9BECD", X"FAE5EA", X"F6F4F5", X"F5F7F6", X"F5F6F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEDF1", X"F9BBCB", X"F4809E", X"F1567E", X"EF426F", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EB416D", X"E73F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"EB416D", X"EF406E", X"EF406D", X"EF4773", X"F26287", X"F28EA8", X"F1C0CD", X"F4EAED", X"F5F7F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFD", X"F9BFCE", X"F36D90", X"EF4672", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EB416D", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E73F6B", X"ED416E", X"EF426F", X"EF426F", X"EF406E", X"EF406E", X"ED4A74", X"ED7594", X"F1C0CD", X"F5F4F4", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FAFAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFE", X"F9B4C6", X"F04F79", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"E9406C", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E8406C", X"ED426E", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"EE3F6D", X"ED527B", X"F4BAC9", X"F9F9F9", X"F9F9F9", X"FBFBFB", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDFE6", X"F15981", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"E8406C", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E8406C", X"EE426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F26B8E", X"FEF0F3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9B7C8", X"EF4572", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"ED426E", X"E8406C", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"EA406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F0517A", X"FCDBE3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9BCCC", X"EF4773", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"EE426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EC416E", X"E73F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"EB416D", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F1547D", X"FCDEE6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBF0", X"F36D90", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426E", X"E9406C", X"E7406C", X"E8406C", X"E9406C", X"E9406C", X"EA406D", X"EA416D", X"EB416D", X"EC416E", X"ED416E", X"ED416E", X"EE426E", X"EE426F", X"EF426F", X"EF426F", X"EB416D", X"E73F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"EC416D", X"EF426F", X"EF416E", X"EF416E", X"F589A5", X"FEF8FA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCD6E0", X"F47999", X"F04874", X"EF406D", X"EF3F6D", X"EF3F6D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"ED3F6C", X"E83D6A", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E63D69", X"E73D6A", X"E73D6A", X"E83D6A", X"E83D6A", X"E93E6B", X"E93E6B", X"E73D6A", X"E63D69", X"E63D69", X"E63D69", X"E63C69", X"E73D69", X"EC406D", X"F04E78", X"F58BA6", X"FDEAEF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF1F4", X"FAC2D1", X"F68FAA", X"F47A9A", X"F36F91", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F26A8E", X"F0698C", X"EA6689", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96688", X"E96689", X"EA6B8D", X"EA7795", X"F096AE", X"FBD0DC", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFD", X"FEF5F7", X"FEF1F4", X"FEF0F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FAEDF1", X"F4E8EB", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EB", X"F4E8EB", X"F4E7EB", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EA", X"F4E7EB", X"F4EDEF", X"F7F5F6", X"FCFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFBFB", X"F5F6F6", X"F5F6F6", X"F5F6F6", X"F5F6F6", X"F5F6F6", X"FAFBFB", X"FCFDFD", X"FBFCFC", X"FAFBFB", X"F9FAFA", X"F9F9F9", X"F8F8F8", X"F7F8F8", X"F7F7F7", X"F6F7F7", X"F6F6F6", X"F5F6F6", X"F5F6F6", X"F5F6F6", X"F5F6F6", X"F5F6F6", X"F8F9F9", X"FDFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FEFEFE", X"FDFDFD", X"FDFDFD", X"FCFCFC", X"FCFCFC", X"FBFBFB", X"FAFAFA", X"FAFAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F6", X"F8F9F9", X"FEFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFE", X"FEF5F8", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF3F6", X"FEF8FA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"FEF0F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF1F4", X"FEF2F5", X"FFFDFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF9FA", X"FEF3F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF4F6", X"FEF3F6", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFA", X"FFFAF0", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFFAF0", X"FEF9EF", X"F9F4EB", X"F5F4F0", X"F5F6F7", X"F5F6F7", X"F5F5F5", X"F5F5F5", X"F5F4F3", X"F5EFE4", X"F5EEE2", X"F9F3E7", X"FFF8EB", X"FFF8EC", X"FFF8EC", X"FFF8EB", X"FFFCF5", X"FEFEFF", X"FBFBFB", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFBF5", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9EF", X"FFFAF2", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFBF3", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9EF", X"FFFAF0", X"FFFDF9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFFAF1", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9EF", X"FFFAF0", X"FFFEFB", X"FFFFFF", X"FFFBF5", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9EF", X"FFF9F0", X"FFFDF9", X"FFFFFF", X"FFFCF5", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9EF", X"FFFBF5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFB", X"FFFAF0", X"FFF9EF", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9F0", X"FFF9EF", X"FFFAF1", X"FFFEFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEDF1", X"F4809E", X"F36F91", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F36E91", X"F79FB6", X"FFFAFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBCEDA", X"F37293", X"F36C8F", X"F36D90", X"F36D90", X"F36D90", X"F36C8F", X"F47D9C", X"FEEFF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8B1C3", X"F36E90", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37092", X"F37495", X"F691AB", X"FBD2DC", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF6E5", X"FFD68E", X"FFBF4F", X"FFBA3E", X"FDB83E", X"FDB83E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFBA3E", X"FEB93E", X"F9B53E", X"F5B33C", X"F5B748", X"F5C97B", X"F5EBD9", X"F7F8F9", X"F6F6F7", X"F5F0E9", X"F5C165", X"F5B035", X"F5B138", X"FAB539", X"FFB839", X"FFB839", X"FFB636", X"FFDB9C", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFEAC6", X"FFCB6E", X"FFBC44", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFBA41", X"FFC661", X"FFE4B5", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFC866", X"FFB93C", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFBB42", X"FFE5B5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF6E6", X"FFC152", X"FFB93D", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93D", X"FFBE4A", X"FFEDCD", X"FFFEFC", X"FFD283", X"FFB83B", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFBA40", X"FFE3B0", X"FFFFFE", X"FFD487", X"FFB83B", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFBC45", X"FFC867", X"FFE9C3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFECCA", X"FFBD49", X"FFB93D", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFB93E", X"FFBA3F", X"FFC256", X"FFDDA0", X"FFFAF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBD0DB", X"F04C76", X"EF3E6C", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3D6B", X"F2678B", X"FEF1F4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04874", X"EF3F6D", X"EF406D", X"EF406D", X"EF406D", X"EF3E6C", X"F15880", X"FDEBF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F696AF", X"EE3C6A", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF3F6D", X"EF406D", X"F1547D", X"F9B7C8", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF1D9", X"FFBC46", X"FFA402", X"FFA200", X"FCA000", X"F69D00", X"F79D00", X"FDA000", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FDA100", X"F89D00", X"F59C00", X"F59C00", X"F59B00", X"F59D00", X"F9B844", X"FEF2DB", X"FAFBFD", X"F5F0E7", X"F5B33E", X"F59B00", X"F59C00", X"F69C00", X"FCA000", X"FFA200", X"FFA100", X"FFD589", X"FFFFFF", X"FFFFFE", X"FFDDA2", X"FFAD1B", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA910", X"FFD386", X"FFFDF9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB532", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA402", X"FFDB9C", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DD", X"FFAB17", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFA70C", X"FFE7BC", X"FFFDFB", X"FFC359", X"FFA000", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFD995", X"FFFEFE", X"FFC45D", X"FFA000", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFAE1F", X"FFE2AF", X"FFFFFF", X"FFFFFF", X"FFE5B8", X"FFA70B", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA506", X"FFC764", X"FFF8EC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9B4C6", X"EF4571", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F1547D", X"FDE1E8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15D83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F15A81", X"FCDEE6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC867", X"FFA200", X"FFA300", X"FBA100", X"F69E00", X"F59D00", X"F59D00", X"F89F00", X"FEA200", X"FFA300", X"FFA300", X"FFA300", X"FCA100", X"F79E00", X"F59D00", X"F59D00", X"F59D00", X"F69D00", X"FAA000", X"FFA200", X"FFCC71", X"FFFEFC", X"F9F4EB", X"F5B440", X"F59C00", X"F59D00", X"F59D00", X"F69E00", X"FDA200", X"FFA301", X"FFD791", X"FFFFFF", X"FFEFD3", X"FFAF21", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA911", X"FFE7BB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFEFB", X"FFC45B", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA402", X"FFD996", X"FFFFFE", X"FFC660", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB532", X"FFF6E5", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA403", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F698B1", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04A75", X"FAC5D3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4471", X"F9B3C5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF6E5", X"FFB024", X"FFA200", X"FEA200", X"F79E00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F99F00", X"FFA300", X"FFA300", X"FCA100", X"F69E00", X"F59D00", X"F59D00", X"F59D00", X"F69E00", X"FBA100", X"FFA300", X"FFA200", X"FFB22B", X"FFF6E7", X"FEF9F1", X"F8B642", X"F59C00", X"F59D00", X"F59D00", X"F89F00", X"FEA200", X"FFA301", X"FFD790", X"FFFFFF", X"FFDA98", X"FFA403", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFCF7A", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFEFB", X"FFC45B", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA402", X"FFD996", X"FFFEFE", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA609", X"FFE2AD", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC152", X"FFFCF5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF7F9", X"F47D9C", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"F8AABE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F7A2B8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DC", X"FFAC19", X"FFA200", X"FFA300", X"FCA100", X"F69D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"FAA000", X"FAA000", X"F69D00", X"F59D00", X"F59D00", X"F59D00", X"F79E00", X"FCA100", X"FFA300", X"FFA300", X"FFA200", X"FFAB17", X"FFF0D7", X"FFFAF2", X"FDBA43", X"F79D00", X"F59D00", X"F99F00", X"FEA200", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD488", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC763", X"FFFDFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFEFB", X"FFC45B", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA402", X"FFD996", X"FFFEFE", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD892", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83B", X"FFF9ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEEDF1", X"F26287", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F68FA9", X"FFFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF416E", X"EF416E", X"EF416E", X"EF416E", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FBA000", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F89F00", X"FDA200", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAB17", X"FFF0D6", X"FFFAF2", X"FFBB43", X"FDA000", X"FBA100", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFEFB", X"FFC45B", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA402", X"FFD996", X"FFFEFE", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD891", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCD9E2", X"F0517A", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F37294", X"FEF4F6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4672", X"F04C77", X"F04C77", X"F04C77", X"F04C77", X"F04C77", X"F04C77", X"EF4572", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FAA000", X"F59D01", X"F5A00A", X"F5A20D", X"F5A20D", X"F5A20D", X"F5A20D", X"F5A20D", X"F9A30C", X"FEA301", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAB17", X"FFF0D6", X"FFFAF2", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA404", X"FFA80D", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA506", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFEFB", X"FFC45B", X"FFA200", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFA403", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFA403", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFA402", X"FFD996", X"FFFEFE", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA506", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80D", X"FFA505", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD892", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA401", X"FFA70C", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA80E", X"FFA608", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FABECD", X"F04873", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F15981", X"FDE7ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F47797", X"FBCBD8", X"FBCEDA", X"FBCEDA", X"FBCEDA", X"FBCFDA", X"FAC9D6", X"F37092", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFDFE", X"FDF1DA", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FEA200", X"F8A30B", X"F5CD88", X"F5DFB8", X"F5DEB6", X"F5DEB6", X"F5DEB6", X"F9E3BB", X"FEDEA5", X"FFAA13", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAB17", X"FFF0D6", X"FFFAF2", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB532", X"FFE3B2", X"FFE8BE", X"FFE7BD", X"FFE7BD", X"FFE7BD", X"FFE7BD", X"FFC154", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC662", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFEFB", X"FFC35A", X"FFA200", X"FFAA12", X"FFB228", X"FFBC45", X"FFCB6E", X"FFDB9D", X"FFC55E", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80D", X"FFD385", X"FFD78F", X"FFC661", X"FFB83B", X"FFAF22", X"FFA70B", X"FFA402", X"FFD996", X"FFFEFE", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC256", X"FFE8BE", X"FFE7BD", X"FFE7BD", X"FFE7BD", X"FFE7BD", X"FFE5B8", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD892", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFAA14", X"FFDFA7", X"FFE8BE", X"FFE7BD", X"FFE7BD", X"FFE7BD", X"FFE8C0", X"FFCC72", X"FFA403", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F7A1B8", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04D77", X"FBCEDA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F58AA6", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"F4819F", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F8F8F8", X"F5F6F8", X"F8EBD4", X"FEAB19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FEA810", X"F7E1BB", X"F5F7FB", X"F5F6F9", X"F5F6F9", X"F5F6F8", X"F8FAFE", X"FEF4E3", X"FFAE1D", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFAB17", X"FFF0D6", X"FFFAF2", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB44", X"FFFBF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCD73", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFE", X"FFE2AF", X"FFDDA0", X"FFE9C3", X"FFF4E1", X"FFFCF7", X"FFFEFD", X"FFFFFF", X"FFD589", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFEAC6", X"FFFFFF", X"FFFEFC", X"FFFBF2", X"FFF1D8", X"FFE6BA", X"FFDA97", X"FFECCA", X"FFFEFB", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD75", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFC55F", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFA301", X"FFD892", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1C", X"FFF6E5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDB9C", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAFB", X"F585A2", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4470", X"F8B2C4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F6F7", X"F5E9D3", X"F8A818", X"FEA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FDE6BD", X"F6F8F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F6", X"F9F6F1", X"FFE3B1", X"FFD282", X"FFC257", X"FFB533", X"FFAD1B", X"FFA505", X"FFAB15", X"FFF0D6", X"FFFAF2", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFECCB", X"FFD790", X"FFC865", X"FFB93D", X"FFB023", X"FFA70C", X"FFA300", X"FFD791", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF1F4", X"F2698D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F696AF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F6F7", X"F6E9D3", X"F9A818", X"FDA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FCFDFF", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F6", X"FAFBFE", X"FFFFFF", X"FFFDFB", X"FFF8ED", X"FFEECF", X"FFE2AF", X"FFD996", X"FFF7EA", X"FFFAF1", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFFBF4", X"FFF2DA", X"FFE6BB", X"FFD997", X"FFEBC7", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCE0E8", X"F1547D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F47999", X"FEF6F8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFBFC", X"FDF0D9", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC5D3", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15E84", X"FDEBF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFF2DC", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8A8BD", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4571", X"EF4370", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04F79", X"FCD5DF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FDA100", X"FCA100", X"FAA000", X"FAA000", X"FCA100", X"FFA810", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFC660", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFD", X"F58DA8", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F2688C", X"F0517A", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4672", X"F9B9CA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCEFD9", X"F8A819", X"F69D00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F9A510", X"FEE7BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCD", X"FFDEA4", X"FFDFA5", X"FFDFA5", X"FFDFA5", X"FFDFA5", X"FFDEA4", X"FFEBC8", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF3F6", X"F37193", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F691AB", X"F37193", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F79EB5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F8F9FA", X"F5E9D3", X"F5A618", X"F59C00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F5A30F", X"FBE4BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FAFAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDE7ED", X"F15980", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4772", X"F9B5C7", X"F58FAA", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F482A0", X"FEF9FA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F8F8F8", X"F6F6F6", X"F5F6F7", X"F5E9D3", X"F5A618", X"F59C00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F5A20F", X"F7E0B9", X"FEFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBCDD9", X"F04D77", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04F79", X"FCD8E1", X"F8AABE", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F2668B", X"FEEFF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FAFAFA", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F6F7", X"F5E9D3", X"F5A618", X"F69D00", X"F89F00", X"F79E00", X"F59D00", X"F59D00", X"F5A20F", X"F6DFB8", X"FEFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8B1C4", X"EF4470", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15E84", X"FEEEF2", X"FAC4D2", X"F04A75", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F0537C", X"FCDEE6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F6F7", X"F6EAD4", X"FAA918", X"FEA100", X"FFA300", X"FCA100", X"F69D00", X"F59D00", X"F5A20F", X"F6E0B9", X"FEFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F696AF", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F47898", X"FEF7F9", X"FCDFE7", X"F0537C", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"F04A75", X"FAC3D1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F4809E", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9FAFB", X"FDF0DA", X"FFAC19", X"FFA200", X"FFA300", X"FBA000", X"F59D00", X"F59D00", X"F5A20F", X"F9E2BB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF6F8", X"F47A99", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F694AD", X"FFFFFF", X"FEF0F3", X"F2668B", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F8A7BC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F698B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F58AA6", X"FFFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAFB", X"F4819F", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9FA", X"FDFDFF", X"FFFFFF", X"FFF3DD", X"FFAC19", X"FFA200", X"FDA200", X"F69E00", X"F59D00", X"F59D00", X"F6A310", X"FCE6BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9ED", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9F", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF4E0", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFB", X"FFC660", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6BA", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDB9B", X"FFA404", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDECF0", X"F15F85", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4370", X"F8AFC2", X"FFFFFF", X"FEF9FA", X"F483A0", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F58BA7", X"FFFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFDFE", X"F9B7C8", X"F586A3", X"F588A4", X"F588A4", X"F26187", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F15C83", X"F586A3", X"F588A4", X"F588A4", X"F588A4", X"F588A4", X"F585A2", X"F15980", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F7F7F7", X"F7F7F7", X"F9F9F9", X"FAFAFA", X"FDFEFF", X"FFEBC8", X"FFC763", X"FFC55E", X"FFC051", X"FFA609", X"FCA100", X"F79E00", X"F59D00", X"F59D00", X"F59D00", X"FAA206", X"FFBC46", X"FFC55F", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC45C", X"FFD282", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFDC9D", X"FFC45B", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC45B", X"FFDB9B", X"FFFEFC", X"FFFFFF", X"FFF8ED", X"FFCC72", X"FFC45D", X"FFC55E", X"FFC257", X"FFAA13", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA402", X"FFB83A", X"FFC55F", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55F", X"FFC052", X"FFA60A", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFCF79", X"FFC45D", X"FFC45C", X"FFB023", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB22B", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC868", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFECCA", X"FFC764", X"FFC55D", X"FFC55F", X"FFBC44", X"FFA505", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA70A", X"FFC153", X"FFC55F", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55F", X"FFB739", X"FFA301", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCD6E0", X"F0507A", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04C77", X"FBCBD7", X"FFFFFF", X"FFFFFF", X"F79EB5", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F36F92", X"FEF3F6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FEF5F8", X"F47697", X"EE3C6A", X"EF3E6C", X"EF3E6C", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF3E6C", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD589", X"FFA100", X"FFA100", X"FFA100", X"FBA000", X"F69E00", X"F59D00", X"F59D00", X"F59D00", X"F99F00", X"FEA200", X"FFA200", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA000", X"FFB636", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFAF2", X"FFBC45", X"FFA000", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA000", X"FFC55E", X"FFFDFA", X"FFFFFF", X"FFECCB", X"FFA910", X"FFA100", X"FFA100", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF0D7", X"FFAB15", X"FFA100", X"FFA100", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA70B", X"FFE7BC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD68E", X"FFA100", X"FFA100", X"FFA100", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA100", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9BACA", X"EF4773", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F1577F", X"FDE4EB", X"FFFFFF", X"FFFFFF", X"F9B9CA", X"EF4672", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F15880", X"FDE6EC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FDEBEF", X"F15D84", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"ED426E", X"EE426F", X"EF426F", X"EF3E6C", X"F7A0B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFB", X"FFC865", X"FFA100", X"FDA200", X"F99F00", X"F59D00", X"F59D00", X"F59D00", X"F59D00", X"F99F00", X"FEA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83A", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFF5E4", X"FFB025", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFDFA6", X"FFA608", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE4B3", X"FFA70C", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA90F", X"FFE7BE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFC969", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB738", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F79EB5", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F36D90", X"FEF2F5", X"FFFFFF", X"FFFFFF", X"FBD5DF", X"F04F79", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04D77", X"FBCDD9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FBD4DE", X"F04F79", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EB416D", X"E73F6B", X"E8406C", X"EB416D", X"ED3F6C", X"F7A2B8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9EF", X"FDB83F", X"FA9F00", X"F69E00", X"F59D00", X"F59D00", X"F59D00", X"F69D00", X"FAA000", X"FEA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83A", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFEAC6", X"FFAA12", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFD282", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD68E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA90F", X"FFE7BE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB42", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB93D", X"FFF9EE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9FA", X"F582A0", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FDEBF0", X"F15D84", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4471", X"F8B2C4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"F9B7C8", X"EF4672", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"EA406D", X"E63F6B", X"E63F6B", X"E63F6B", X"E63E6B", X"E7436E", X"F3B7C7", X"FCFFFE", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFCFD", X"F8EDD8", X"F6A81E", X"F59C00", X"F59D00", X"F59D00", X"F59D00", X"F69E00", X"FBA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83A", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFDDA1", X"FFA506", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFB", X"FFFDF9", X"FFC55D", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFC96A", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA90F", X"FFE7BE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF4E0", X"FFAF20", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC55F", X"FFFDF9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEEFF3", X"F2668A", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F7A3B9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF5F7", X"F47797", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F697B0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"F79BB3", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"E9406C", X"E63F6B", X"E63F6B", X"E63F6B", X"E63E6B", X"E63C69", X"EA6E8F", X"F3E4E8", X"F6F7F6", X"F7F7F7", X"FBFBFB", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFBFD", X"F5DEB4", X"F5A20E", X"F59D00", X"F59D00", X"F59D00", X"F89F00", X"FDA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83A", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFD07D", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFEFB", X"FFF9ED", X"FFB737", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBC44", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA90F", X"FFE7BE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE8BF", X"FFA910", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAB15", X"FFE5B8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCDEE6", X"F0527C", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"F04974", X"FAC1D0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F694AD", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F47C9B", X"FEF7F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDEDF1", X"FEF9FA", X"F47D9C", X"EF3D6B", X"EF406D", X"EF406D", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"ED416E", X"E73E6B", X"E63D69", X"E63D69", X"E63D69", X"E6456F", X"EA7191", X"F2D3DB", X"F5F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFFFF", X"F9D390", X"F59D00", X"F59C00", X"F79D00", X"FBA000", X"FEA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFB737", X"FFF8ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFCF6", X"FFC255", X"FFA100", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFEFC", X"FFF1D8", X"FFAB17", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF4E1", X"FFAE1F", X"FFA100", X"FFA200", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA80D", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD996", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA301", X"FFB126", X"FFDC9E", X"FFFEFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F9B4C6", X"F79EB5", X"F7A0B7", X"F585A2", X"EF4773", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4874", X"F589A5", X"F7A0B7", X"F79FB6", X"F79FB6", X"F7A1B7", X"F37294", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F26086", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDEDF1", X"FFFAFB", X"F9B7C8", X"F7A1B7", X"F7A2B8", X"F7A2B8", X"F7A2B8", X"F36D90", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"F04E78", X"EF4571", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EE426F", X"EC7291", X"ED9DB2", X"ED9BB0", X"EEA1B5", X"F3C0CD", X"F6E9EC", X"F5F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"FBFBFB", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEE7BE", X"FACD7E", X"FBCF81", X"FED182", X"FFCB6F", X"FFA80D", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA608", X"FFC661", X"FFD283", X"FFD281", X"FFD281", X"FFD281", X"FFD180", X"FFDC9E", X"FFFCF6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFCF7", X"FFDDA0", X"FFD180", X"FFD281", X"FFB839", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC662", X"FFFEFB", X"FFF4E2", X"FFD589", X"FFD180", X"FFD281", X"FFD282", X"FFCE77", X"FFAD1B", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA403", X"FFC050", X"FFD283", X"FFD281", X"FFD281", X"FFD281", X"FFD282", X"FFCB70", X"FFA80D", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF6E7", X"FFD58B", X"FFD180", X"FFD281", X"FFD17E", X"FFB430", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83B", X"FFD282", X"FFD281", X"FFD281", X"FFD281", X"FFD180", X"FFD489", X"FFF3DF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE9C1", X"FFD17F", X"FFD281", X"FFD281", X"FFD283", X"FFC55E", X"FFA607", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFA910", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAF22", X"FFCF7B", X"FFD281", X"FFD283", X"FFDC9D", X"FFF1D8", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDE8EE", X"F15A81", X"EF406E", X"EF426F", X"EF416F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F0507A", X"FCD7E0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F47898", X"F2688C", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"ED7494", X"F4EAED", X"F5F6F6", X"F5F6F6", X"FAFDFC", X"FEFFFF", X"FBFBFB", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"F9F9F9", X"FDFDFD", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DC", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC72", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EC", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFA", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAC1A", X"FFC55E", X"FFA402", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAB17", X"FFEAC4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBD0DB", X"F04E78", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4773", X"F9BACB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F58BA6", X"F8ACBF", X"EF4571", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"EB4772", X"F0B6C5", X"F5F7F7", X"F5F5F5", X"F8F8F8", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"FDFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DC", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EC", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFA", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD73", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAE1E", X"FFE5B6", X"FFAF21", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC660", X"FFFDF8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F8B4C6", X"EF4571", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F79EB5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F58BA6", X"FDE5EC", X"F2668B", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EC3F6C", X"EA6E8E", X"F4E7EB", X"F5F6F6", X"F6F6F6", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1C", X"FFF4DF", X"FFCC72", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFAA13", X"FFE7BE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F698B0", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F4819F", X"FEF8FA", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F58AA6", X"FFFCFC", X"F8A7BC", X"EF4370", X"EF426F", X"EF426F", X"EF426F", X"EE416E", X"E7456F", X"EFB1C2", X"F5F7F6", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFA", X"FFD996", X"FFCD75", X"FFDC9E", X"FFE9C4", X"FFF3DD", X"FFF9EE", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF6E4", X"FFECCC", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC45A", X"FFFCF6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF7F9", X"F47C9B", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F26589", X"FEEFF3", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F589A5", X"FFFDFD", X"FDE4EB", X"F15F85", X"EF406E", X"EF426F", X"EF426F", X"EE426F", X"E83E6B", X"EA6A8C", X"F4E6E9", X"F5F6F6", X"FAFAFA", X"FEFEFE", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"F8F8F8", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB43", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC71", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD74", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCF8", X"FFC358", X"FFA100", X"FFA505", X"FFA70D", X"FFAF22", X"FFBA41", X"FFC660", X"FFEAC4", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFEFC", X"FFC866", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE6B9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDECF1", X"F15E85", X"EF3E6C", X"EF406D", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F0527B", X"FCDBE4", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6C", X"EF426F", X"EF426F", X"EC416E", X"EB416D", X"EF3F6D", X"F589A5", X"FFFBFC", X"FFFFFF", X"F79EB5", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EA406C", X"E6436E", X"EFADBE", X"F5F7F6", X"F8F8F8", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBB44", X"FFFBF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCC73", X"FFA100", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFCD75", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFB", X"FFC45C", X"FFA200", X"FFA300", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFD790", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFE9C1", X"FFAA14", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC255", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF0F4", X"F8A8BC", X"F79EB5", X"F79DB4", X"F2658A", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F26288", X"F79CB3", X"F79FB6", X"F79FB6", X"F79FB6", X"F79FB6", X"F79FB6", X"F79FB6", X"F694AE", X"F04D77", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416F", X"F04874", X"FABFCE", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EF3F6D", X"EF426F", X"EB416D", X"E63F6B", X"E73F6B", X"EB3E6B", X"F589A5", X"FFFBFC", X"FFFFFF", X"FCDFE6", X"F15A81", X"EF416E", X"EF426F", X"EF426F", X"EB416D", X"E63D69", X"E96789", X"F4E4E8", X"F5F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAF22", X"FFCF7A", X"FFD282", X"FFD282", X"FFD282", X"FFD282", X"FFD282", X"FFB83A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC662", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EC", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC560", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB83B", X"FFD282", X"FFD282", X"FFD282", X"FFD282", X"FFD282", X"FFD17E", X"FFB42E", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD892", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFCF7", X"FFC359", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE4B5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF5F8", X"F37898", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F697AF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF1F4", X"F2698D", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F7A4B9", X"FFFFFF", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697B0", X"EE3E6C", X"E9406D", X"E63F6B", X"E63F6B", X"E63F6B", X"E73C69", X"F288A4", X"FFFBFC", X"FFFFFF", X"FFFDFE", X"F695AE", X"EF416E", X"EF426F", X"EF426F", X"ED416E", X"E73F6B", X"E6426D", X"EFAABC", X"F5F6F6", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD892", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFE4B5", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC051", X"FFFBF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDEBF0", X"F15D84", X"EF406E", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF4470", X"F9B1C4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAFB", X"F585A2", X"EF3F6D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF3F6D", X"F588A5", X"FFFBFC", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F597AF", X"E83D6A", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63C69", X"ED85A1", X"FDF9FA", X"FFFFFF", X"FFFFFF", X"FCD7E0", X"F0547C", X"EF416E", X"EF426F", X"EE426F", X"E8406C", X"E63D69", X"E96688", X"F3E3E7", X"F6F7F6", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC661", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD891", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFAF2", X"FFBE4C", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80D", X"FFE3B2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBD5DF", X"F04F79", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04D77", X"FBCDD9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F7A0B6", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F36D90", X"FEF2F5", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F496AE", X"E63C69", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63C69", X"EB849F", X"F7F4F5", X"FEFEFE", X"FFFFFF", X"FFFBFC", X"F58BA6", X"EF406D", X"EF426F", X"EF426F", X"E9406C", X"E63F6B", X"E6426D", X"EEA8BB", X"F8F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFD489", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA100", X"FFC764", X"FFFEFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA402", X"FFD894", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA8", X"FFA609", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFC04F", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9BACA", X"EF4672", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F1587F", X"FDE6EC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9BBCB", X"EF4773", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F1577F", X"FDE4EB", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15C83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F597AF", X"E73C69", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63C69", X"EC849F", X"F5F1F2", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FBCEDA", X"F04F79", X"EF416E", X"EF426F", X"EB416D", X"E63F6B", X"E63D69", X"E96487", X"F5E4E8", X"FEFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD790", X"FFFFFF", X"FFDEA3", X"FFA506", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFD17F", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA70B", X"FFE4B4", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EC", X"FFBA3F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA70C", X"FFE3B0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F79FB6", X"EF406D", X"EF426F", X"EF426F", X"EF426F", X"EF426F", X"EF406D", X"F36F91", X"FEF3F6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCD7E0", X"F0507A", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF416E", X"F04C77", X"FBCBD7", X"FFFFFF", X"FAC4D2", X"F04A75", X"EF416E", X"EF426F", X"EF426F", X"EF426F", X"EF406E", X"F15D83", X"FDECF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F697AF", X"E83C69", X"E63F6B", X"E63F6B", X"E63F6B", X"E63F6B", X"E63C69", X"EC849F", X"F5F1F2", X"F5F6F5", X"FAFAFA", X"FFFFFF", X"FEF7F9", X"F47F9E", X"EF406D", X"EF426F", X"EC416E", X"E63F6B", X"E63F6B", X"E6426D", X"EFA8BA", X"FDFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAC19", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA910", X"FFE8BF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBB43", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA301", X"FFD791", X"FFFFFF", X"FFF4E1", X"FFB636", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAE20", X"FFECCB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB635", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA505", X"FFDC9E", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFAC1A", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA80F", X"FFE7BD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD487", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA911", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55F", X"FFA200", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFB93D", X"FFF7E9", X"FFFFFF", X"FFE6B9", X"FFA80E", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFAD1B", X"FFF5E2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDA9A", X"FFA505", X"FFA300", X"FFA300", X"FFA300", X"FFA300", X"FFA200", X"FFBF4D", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9FA", X"F4819F", X"EF3D6B", X"EF406D", X"EF406D", X"EF406D", X"EF406D", X"EF3D6B", X"F58AA6", X"FFFCFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDECF0", X"F15D84", X"EF3E6C", X"EF406D", X"EF406D", X"EF406D", X"EF3F6D", X"EF416E", X"F8AEC1", X"FFFFFF", X"FAC3D2", X"F04873", X"EF3F6D", X"EF406D", X"EF406D", X"EF406D", X"EF3E6C", X"F1577F", X"FDEBF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F696AF", X"E93B68", X"E63D69", X"E63D69", X"E63D6A", X"E93E6B", X"E63A67", X"EB829E", X"F5F1F2", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FAC3D1", X"F04974", X"EF3F6D", X"ED3F6D", X"E73D6A", X"E63D69", X"E63B68", X"E96185", X"FAE6EB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFAB16", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFA80D", X"FFE7BE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBA41", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFD68C", X"FFFFFF", X"FFFFFF", X"FFE7BC", X"FFB42F", X"FFA300", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFAF21", X"FFDFA6", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFB532", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA402", X"FFDB9C", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DD", X"FFAB17", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFA70C", X"FFE7BC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD385", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFA80E", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFC55E", X"FFA000", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA200", X"FFA402", X"FFB635", X"FFE9C2", X"FFFFFF", X"FFFFFF", X"FFE5B8", X"FFA70B", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFAC18", X"FFF4E1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF6E5", X"FFB533", X"FFA100", X"FFA200", X"FFA200", X"FFA200", X"FFA100", X"FFA608", X"FFE1AB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF7F9", X"F7A4B9", X"F586A3", X"F587A4", X"F587A4", X"F587A4", X"F587A4", X"F586A3", X"FAC3D1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEF8FA", X"F7A6BB", X"F586A3", X"F587A4", X"F587A4", X"F587A4", X"F587A4", X"F585A3", X"FAC0CF", X"FFFFFF", X"FBD3DE", X"F58CA7", X"F589A5", X"F58AA5", X"F58AA5", X"F58AA5", X"F589A5", X"F696AF", X"FEF2F5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FABDCD", X"F183A0", X"EB829E", X"EB829E", X"EB829E", X"F185A1", X"F084A0", X"EFAEBF", X"F5F3F3", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFDFD", X"FEF4F7", X"F79EB5", X"F586A3", X"F487A4", X"EE83A0", X"EB829E", X"EC829E", X"F189A4", X"FBD6E0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF7E8", X"FFCB6E", X"FFC55D", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC868", X"FFF0D7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBF3", X"FFD282", X"FFC55F", X"FFC661", X"FFC661", X"FFC661", X"FFC661", X"FFC55E", X"FFE3B1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFD791", X"FFC866", X"FFC55D", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC762", X"FFD488", X"FFEECF", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBF3", X"FFD17F", X"FFC45C", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC661", X"FFE9C1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFCB6F", X"FFC45D", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC867", X"FFF0D5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE4B3", X"FFC45C", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC969", X"FFF1D9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFDB9A", X"FFC45B", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55D", X"FFC968", X"FFDA99", X"FFF3DE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEFD3", X"FFC867", X"FFC55D", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC45D", X"FFCB6F", X"FFF9ED", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A8", X"FFC45C", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC55E", X"FFC45B", X"FFDB9C", X"FFFEFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBFC", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFBFC", X"FFFDFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCFD", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFAFC", X"FFFCFD", X"FFFFFF", X"FFFCFD", X"FFFBFC", X"FFFBFC", X"FFFBFC", X"FFFBFC", X"FFFBFC", X"FFFBFC", X"FFFBFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFD", X"FCF8F9", X"F5F1F2", X"F5F1F2", X"F4F1F2", X"F9F5F6", X"FEFAFB", X"F9F6F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFCFD", X"FFFAFC", X"FFFAFC", X"F9F5F6", X"F6F2F3", X"FBF7F8", X"FEFAFB", X"FFFCFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFDFA", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFDF9", X"FFFDFA", X"FFFDFA", X"FFFDFA", X"FFFDFA", X"FFFDFA", X"FFFDF9", X"FFFEFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFB", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFA", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFDFA", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFB", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFEFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDFA", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFD", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDF9", X"FFFDFA", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F6F7F7", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FCFDFD", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FEFEFE", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FBFBFB", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FCFCFC", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFD", X"F7F8FA", X"F5F6F8", X"F5F6F9", X"F5F6F9", X"F5F6F9", X"F5F6F9", X"F5F6F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"FBFBFB", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFFFF", X"FDFEFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF7E8", X"FFDD9F", X"FFF8EC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"F9EBD1", X"F5CE88", X"F5CC82", X"F5CC82", X"F5CC82", X"F5CC82", X"F5CB81", X"F5E1BF", X"F5F6F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FCFCFC", X"FEFEFE", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFE", X"FFFFFF", X"FFE7BC", X"FFD385", X"FFD487", X"FFD488", X"FFD58A", X"FFD489", X"FFD487", X"FFD487", X"FFD78F", X"FFF5E3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE4B5", X"FFDA98", X"FFFCF8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFECC9", X"FFD282", X"FFCB6E", X"FFD17F", X"FFE4B4", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF1D8", X"FFD68E", X"FFD487", X"FFD487", X"FFD487", X"FFD487", X"FFD58B", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEBC8", X"FFE1AB", X"FFFDF8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDF9", X"FFECCC", X"FFD893", X"FFCD75", X"FFCE76", X"FFD58C", X"FFE9C3", X"FFFCF6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF1D8", X"FFDFA6", X"FFFCF5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCD", X"FFE2AE", X"FFFDF9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBF5", X"FFDC9D", X"FFD486", X"FFD487", X"FFD488", X"FFD58A", X"FFD488", X"FFD487", X"FFD386", X"FFDEA4", X"FFFCF7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCD", X"FFB42E", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEDDA4", X"F7A81C", X"F5BA50", X"F5BC57", X"F5BC56", X"F5BC56", X"F6BC55", X"F8DDAC", X"F7F8F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFDEA2", X"FFC257", X"FFC45A", X"FFC255", X"FFAD1B", X"FFB635", X"FFC45B", X"FFC359", X"FFC765", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD384", X"FFC051", X"FFFCF6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDEA5", X"FFB22A", X"FFBD47", X"FFC867", X"FFC662", X"FFBC45", X"FFE4B4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A9", X"FFAD1C", X"FFC152", X"FFC45A", X"FFC45A", X"FFC359", X"FFC55F", X"FFEBC6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF4F", X"FFFBF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBF4", X"FFD07C", X"FFB229", X"FFBD48", X"FFC662", X"FFC867", X"FFC256", X"FFBB43", X"FFEAC5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0AA", X"FFB93C", X"FFF7EA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD792", X"FFBF4E", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFCE78", X"FFC358", X"FFC45B", X"FFBD48", X"FFA911", X"FFBF4C", X"FFC45B", X"FFC358", X"FFD281", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDDA2", X"FDB83E", X"F6EDDD", X"F5F3EF", X"F5F2ED", X"F5F2ED", X"F5F2ED", X"F9F8F5", X"FDFDFD", X"FBFBFB", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FAFAFA", X"FFFFFF", X"FFFDFB", X"FFFCF7", X"FFFDF8", X"FFF7EA", X"FFBD48", X"FFD790", X"FFFEFB", X"FFFCF7", X"FFFCF8", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD997", X"FFC96A", X"FFFEFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF7E8", X"FFB83A", X"FFD489", X"FFFBF3", X"FFFEFC", X"FFFDFA", X"FFF5E4", X"FFF6E7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA6", X"FFB83C", X"FFF5E3", X"FFFDF9", X"FFFCF7", X"FFFCF7", X"FFFCF7", X"FFFEFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF4F", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDB9A", X"FFB32C", X"FFE2AE", X"FFFAF2", X"FFFDFB", X"FFFEFC", X"FFFCF6", X"FFF5E3", X"FFF9EF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A9", X"FFB83B", X"FFF7EA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD791", X"FFBE4D", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFDF9", X"FFFCF7", X"FFFDFA", X"FFEAC6", X"FFB32C", X"FFEFD2", X"FFFDF9", X"FFFCF7", X"FFFDF9", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDDA1", X"FFBA41", X"FCF5EA", X"F6F6F8", X"F5F5F6", X"F5F5F6", X"F5F5F6", X"F5F5F6", X"FAFAFA", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF2", X"FFBE4B", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE7BC", X"FFDFA8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF1DA", X"FFB229", X"FFEAC4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA6", X"FFB93E", X"FFF8EB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF50", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBD47", X"FFD386", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0AA", X"FFB83B", X"FFF7EA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD791", X"FFBF4D", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32E", X"FFF1D9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDDA1", X"FFBB42", X"FFFAF0", X"FBFDFF", X"F5F7FA", X"F5F6F9", X"F5F6F8", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBE4A", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFB", X"FFFDFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF0", X"FFBF4D", X"FFBF4E", X"FFEBC8", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA6", X"FFB93E", X"FFF9EF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF50", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF2DB", X"FFB42F", X"FFEAC5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A9", X"FFB93C", X"FFF9EE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD894", X"FFBF4D", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F8F8F8", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFDEA3", X"FFAF20", X"FFC867", X"FFCB70", X"FAC76D", X"F5C36A", X"F5D191", X"F5F2ED", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F9F9F9", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBE4A", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEFD3", X"FFC45C", X"FFB531", X"FFBD49", X"FFCF7B", X"FFEFD3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA8", X"FFAE20", X"FFC867", X"FFCC71", X"FFCB70", X"FFCB6E", X"FFE0A8", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF50", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFECCB", X"FFB32D", X"FFF1D9", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFCF7A", X"FFCB6F", X"FFCB70", X"FFE2AF", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE1AB", X"FFAE20", X"FFC866", X"FFCC71", X"FFCB70", X"FFCB70", X"FFCC72", X"FFB93E", X"FFBE4C", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFDEA3", X"FFAE20", X"FFC763", X"FFCA6C", X"FEC96B", X"F8C468", X"F5D08E", X"F5F2ED", X"F5F5F6", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBE4A", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCF7", X"FFEECF", X"FFD68D", X"FFBB42", X"FFB531", X"FFE5B8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A8", X"FFAE1F", X"FFC662", X"FFCA6C", X"FFCA6B", X"FFC969", X"FFDFA5", X"FFFEFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF50", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCE", X"FFB32E", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFF3DD", X"FFCD76", X"FFCA6B", X"FFB229", X"FFC867", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE1AB", X"FFAE1F", X"FFC662", X"FFCA6C", X"FFCA6B", X"FFCA6B", X"FFCA6D", X"FFB83B", X"FFBE4C", X"FFFAF3", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D6", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"FCFCFC", X"FFFFFF", X"FFDDA2", X"FFBA40", X"FFF8EB", X"FFFFFF", X"FFFEFD", X"FEFDFC", X"F7F7F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBE4A", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF9EF", X"FFCB6F", X"FFBE4B", X"FFFAF1", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA6", X"FFB93D", X"FFF7E9", X"FFFFFF", X"FFFEFD", X"FFFEFD", X"FFFFFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF50", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DF", X"FFB430", X"FFE8C0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFFFFE", X"FFCA6D", X"FFC868", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0AA", X"FFB83B", X"FFF7E8", X"FFFFFF", X"FFFEFD", X"FFFEFD", X"FFFFFF", X"FFD790", X"FFBF4D", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF0D7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDDA1", X"FFBA41", X"FFF9EE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFE", X"F6F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBE4A", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE5B8", X"FFB42F", X"FFF5E4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA6", X"FFB93E", X"FFF8EB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF50", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFBF3", X"FFBF4D", X"FFD07D", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFCB6F", X"FFC868", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0AA", X"FFB83B", X"FFF7EA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD792", X"FFBF4D", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32D", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCC", X"FFB32B", X"FFECC9", X"FFFAF2", X"FFFAF0", X"FFFAF0", X"FFFAF0", X"FFFCF7", X"FFFFFF", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDDA2", X"FFB93D", X"FFF3DE", X"FFFAF1", X"FFFAF0", X"FFFAF0", X"FFFAF0", X"FCF9F5", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBE4A", X"FFD995", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF2", X"FFE6BB", X"FFF5E4", X"FFFBF4", X"FFFCF7", X"FFF6E6", X"FFCA6C", X"FFBC44", X"FFF9EF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDFA6", X"FFB93D", X"FFF8EB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFBF4F", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFDEA4", X"FFB22A", X"FFDFA7", X"FFF9EE", X"FFFDF9", X"FFFCF6", X"FFF8EB", X"FFC55F", X"FFC866", X"FFFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A9", X"FFB83B", X"FFF7E9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD791", X"FFBE4C", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFECCC", X"FFB32D", X"FFF1D8", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEECF", X"FFAF20", X"FFBA3F", X"FFBF4C", X"FFBE4C", X"FFBE4C", X"FFBD48", X"FFDC9F", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FDFDFD", X"FBFCFF", X"F9DAA2", X"F9A91B", X"FBBA46", X"FEBE4C", X"FFBE4C", X"FFBE4B", X"FFBE4A", X"FFE0AA", X"FBFCFE", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFAF1", X"FFBF4E", X"FFDA97", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EB", X"FFBE4A", X"FFB533", X"FFBE4B", X"FFC052", X"FFB533", X"FFB42E", X"FFE5B7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE0A8", X"FFBA41", X"FFF8EB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD58B", X"FFC050", X"FFFBF4", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFCF7", X"FFD58B", X"FFB530", X"FFBD47", X"FFC45C", X"FFC256", X"FFBC46", X"FFB42E", X"FFDA98", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFE1AB", X"FFBA3F", X"FFF7EA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFD893", X"FFC050", X"FFFAF2", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCD", X"FFB531", X"FFF1D9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8ED", X"FFDFA7", X"FFDB9C", X"FFDB9C", X"FFDB9C", X"FFDB9C", X"FFDB9A", X"FFECCA", X"FCFCFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F8F8F8", X"F6F6F6", X"F5F6F6", X"F5E9D4", X"F5D59B", X"F5D396", X"F7D496", X"FDDA9A", X"FFDB9C", X"FFDB9B", X"FFEED0", X"FFFFFF", X"F9F9F9", X"F5F5F5", X"F8F8F8", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFDFA", X"FFE7BB", X"FFF1D7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFE", X"FFF3DE", X"FFDEA3", X"FFD386", X"FFD283", X"FFD996", X"FFF0D5", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DE", X"FFE5B6", X"FFFCF7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFEDCE", X"FFE5B6", X"FFFDF9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFEFC", X"FFF1D9", X"FFDFA6", X"FFD58B", X"FFD893", X"FFE2AF", X"FFF1DA", X"FFFDF9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF3DF", X"FFE5B6", X"FFFCF7", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF0D6", X"FFE7BC", X"FFFDFA", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFF8EC", X"FFE3B0", X"FFFAF0", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFFFF", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F6F6", X"F5F6F9", X"F5F6F9", X"F5F6F9", X"F9FAFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FBFBFB", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FBFBFB", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FEFEFE", X"FCFCFC", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FAFAFA", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F8F8F8", X"F8F8F8", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FDFDFD", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FAFAFA", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F9F9F9", X"F8F8F8", X"F9F9F9", X"FAFAFA", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"FAFAFA", X"F9F9F9", X"F8F8F8", X"F8F8F8", X"FAFAFA", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"F9F9F9", X"FDFDFD", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"FAFAFA", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F6F6F6", X"F5F5F5", X"F6F6F6", X"FAFAFA", X"FBFBFB", X"FCFCFC", X"FCFCFC", X"FAFAFA", X"F7F7F7", X"F5F5F5", X"F7F7F7", X"FCFCFC", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FDFDFD", X"FAFAFA", X"F7F7F7", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F9F9F9", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF"),
        (X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FEFEFE", X"F7F7F7", X"F5F5F5", X"F8F8F8", X"FDFDFD", X"FDFDFD", X"F9F9F9", X"F8F8F8", X"FEFEFE", X"FFFFFF", X"FDFDFD", X"F8F8F8", X"F5F5F5", X"F7F7F7", X"FEFEFE", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FCFCFC", X"F9F9F9", X"F6F6F6", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F5F5F5", X"F6F6F6", X"FBFBFB", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF", X"FFFFFF")
    );

end endgame_pkg;
